##==========================================================================
##
##      hal_cortexm_kinetis_twr_k60n512_fxm.cdl
##
##      Cortex-M Freescale TWR-K60N512 + TWR-FXM platform HAL configuration
##
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2011 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
##==========================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):    Ilija Kocho <ilijak@siva.com.mk>
## Date:         2011-09-26
##
######DESCRIPTIONEND####
##
##==========================================================================

cdl_package CYGPKG_HAL_CORTEXM_KINETIS_TWR_K60N512_FXM {
    display       "Freescale Kinetis TWR-K60N512-FXM Platform"
    parent        CYGPKG_HAL_CORTEXM_KINETIS
    define_header hal_cortexm_kinetis_twr_k60n512_fxm.h
    include_dir   cyg/hal
    hardware
    requires      { CYGHWR_HAL_CORTEXM_SYSTICK_CLK_SOURCE == "INTERNAL" }

    implements    CYGINT_HAL_CORTEXM_KINETIS_RTC
    implements    CYGINT_IO_FREESCALE_I2C0
    implements    CYGINT_IO_SERIAL_FREESCALE_UART4
    implements    CYGINT_HAL_FREESCALE_UART4

    description   "
    The Freescale TWR K60N512 FXM Platform package provides the support
    needed to run eCos on the TWR K60N512 development system equipped
    with TWR-FXM external memory board. This package
    can also be used for other boards that employ a controller from Kinetis
    families."

    compile       twr_k60n512_fxm_misc.c

    requires      { is_active(CYGPKG_DEVS_ETH_PHY) implies
        (1 == CYGHWR_DEVS_ETH_PHY_KSZ8041) }
    requires      { is_active(CYGPKG_HAL_FREESCALE_EDMA) implies
        (CYGNUM_HAL_FREESCALE_EDMA_CHAN_NUM == 16) }

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_cortexm_kinetis_twr_k60n512_fxm.h>"
        puts $::cdl_header "#define HAL_PLATFORM_CPU    \"Cortex-M4\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Freescale TWR-K60N512-FXM\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
    }

    cdl_component CYG_HAL_STARTUP_ENV {
        display "Startup type"
        flavor data
        no_define
        calculated {
            !CYG_HAL_STARTUP_PLF ? CYG_HAL_STARTUP :
            ((CYG_HAL_STARTUP_PLF == "ByVariant") ?
            (CYG_HAL_STARTUP . "(Variant)") :
            (CYG_HAL_STARTUP . "(Platform)"))
        }
        description "
            Startup type configuration defines the system memory layout.
            Startup type  can be defined by the variant (CYG_HAL_STARTUP_VAR)
            or a platform (CYG_HAL_STARTUP_PLF). If CYG_HAL_STARTUP_PLF
            is defined and not equal to 'ByVariant' then it shall
            override CYG_HAL_STARTUP_VAR."
    }

    cdl_option CYG_HAL_STARTUP_PLF {
        display       "By platform"
        flavor        data
        parent        CYG_HAL_STARTUP_ENV
        default_value { "ROM" }
        legal_values  { "ByVariant" "ROM" "RAM" }
        requires      { CYG_HAL_STARTUP_PLF != "ByVariant" implies
                        CYGPKG_HAL_CORTEXM_KINETIS_FBRAM == 1 }

        description   "
            Startup tupes provided by the platform, in addition to variant
            startup types.
            If 'ByVariant' is selected, then startup type shall be selected from
            the variant (CYG_HAL_STARTUP_VAR). Platform's 'ROM' startup builds
            application similar to Variant's 'ROM' but using external RAM (FlexBus).
            'RAM' startup builds application intended for loading by RedBoot into
            external RAM."
    }

    cdl_component CYGHWR_MEMORY_LAYOUT_PLF {
        display "Memory layout by platform"
        flavor data
        no_define
        active_if { CYG_HAL_STARTUP_PLF != "ByVariant" }
        implements CYGINT_HAL_CORTEXM_KINETIS_FBRAM
        parent  CYGHWR_MEMORY_LAYOUT
        calculated {
            (CYG_HAL_STARTUP_PLF == "ByVariant" ) ? "by variant" :
            (CYG_HAL_STARTUP == "RAM") ? "kinetis_"
            . CYGHWR_HAL_CORTEXM_KINETIS_OC_MEM_LAYOUT  . "_extram_ram" :
            (CYG_HAL_STARTUP == "ROM") ? "kinetis_"
            . CYGHWR_HAL_CORTEXM_KINETIS_OC_MEM_LAYOUT  . "_extram_rom" :
            "Error!" }
        description "Combination of 'Startup type' and 'Kinetis member in use'
        produces the memory layout."

        cdl_option CYGHWR_MEMORY_RAM_RESERVED {
            display "Reserved RAM space \[Bytes\]"
            flavor  data
            legal_values 0 to 0x40000
            default_value 0x20000
        }
    }

    cdl_option CYGHWR_HAL_CORTEXM_KINETIS_PLF_XTAL_OR_OSC_FREQ {
        display "Platform Clock Frequency"
        flavor data
        parent CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT
        default_value 50000000
        legal_values { 25000000 50000000 }
    }

    cdl_option CYGHWR_HAL_CORTEXM_KINETIS_PLF_OSC_CAP {
        display "Platform requred XTAL || C \[pF\]"
        flavor bool
        default_value { CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT_IS == "XTAL" }
        parent CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT
        active_if { CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT_IS == "XTAL" }
        requires { CYGHWR_HAL_CORTEXM_KINETIS_OSC_CAP == 20 }
    }

    cdl_option CYGHWR_HAL_CORTEXM_KINETIS_PLF_RTC {
        display "Platform requred RTC XTAL || C \[pF\]"
        flavor bool
        default_value 1
        parent CYGHWR_HAL_CORTEXM_KINETIS_RTC
        requires { CYGHWR_HAL_CORTEXM_KINETIS_RTC_OSC_CAP == 20 }
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        legal_values 0 to 2
        default_value   1
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
        The TWR board has one serial port fitted to RS232 connector. This option
        chooses which port will be used to connect to a host
        running GDB."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
        display          "Diagnostic serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
        The TWR has one serial port fitted to RS232 connector. This option
        chooses which port will be used for diagnostic output."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Console serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 38400
        description   "
        This option controls the default baud rate used for the
        console connection.
        Note: this should match the value chosen for the GDB port if the
        diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 38400
        description   "
        This option controls the default baud rate used for the
        GDB connection.
        Note: this should match the value chosen for the console port if the
        console and GDB port are the same."
    }

    cdl_component CYGHWR_DEVS_DISK_MMC_FREESCALE_DSPI_BUS {
        display "MMC Disk SPI bus"
        flavor data
        parent CYGPKG_DEVS_DISK_MMC_FREESCALE_DSPI
        calculated 1

        requires CYGHWR_DEVS_SPI_FREESCALE_DSPI1 == 1
        implements CYGINT_DEVS_SPI_FREESCALE_DSPI1
        implements CYGINT_FREESCALE_DSPI1_HAS_MASS

        cdl_option CYGHWR_DEVS_DISK_MMC_FREESCALE_DSPI_CS {
            display "Device number (CS)"
            flavor data
            calculated 0
            implements CYGINT_FREESCALE_DSPI1_CS0
        }
    }

    cdl_option CYGNUM_DEVS_FLASH_SPI_SST25XX_DEV0_MAP_ADDR {
        display "SST25XX Flash Mapping Address"
        flavor data
        parent CYGHWR_DEVS_FLASH_SPI_SST25XX_DEV0
        default_value 0xD0000000
    }
    cdl_component CYGHWR_DEVS_FLASH_SST25XX_DEV0_SPI_BUS {
        display "SST25xx SPI bus"
        flavor data
        parent CYGHWR_DEVS_FLASH_SPI_SST25XX_DEV0
        calculated 1

        requires CYGHWR_DEVS_SPI_FREESCALE_DSPI1 == 1
        implements CYGINT_DEVS_SPI_FREESCALE_DSPI1

        cdl_option CYGHWR_DEVS_FLASH_SST25XX_DEV0_SPI_CS {
            display "Device number (CS)"
            flavor data
            calculated 1
            implements CYGINT_FREESCALE_DSPI1_CS1
        }
    }

    cdl_component CYGHWR_HAL_DEVS_IRQ_PRIO_SCHEME {
        display "Interrupt priority scheme"
        flavor none
        description "Consolidated interrupt priority scheme setting."
    }

    cdl_component CYGPKG_HAL_EXTRN_MEMORY {
        display "External memory devices"
        parent CYGPKG_HAL_CORTEXM_KINETIS_FLEXBUS
        flavor none
        active_if {
            CYGHWR_HAL_KINETIS_FB_CS0 || CYGHWR_HAL_KINETIS_FB_CS1 ||
            CYGHWR_HAL_KINETIS_FB_CS2 || CYGHWR_HAL_KINETIS_FB_CS3 ||
            CYGHWR_HAL_KINETIS_FB_CS4 || CYGHWR_HAL_KINETIS_FB_CS5
        }
        description "
        This is a container for  memory devices attached to
        external bus such as RAM, FLASH, etc."
    }
# FlexBus Implementation
    implements CYGINT_HAL_CORTEXM_KINETIS_FLEXBUS
    implements CYGINT_HAL_EXTRN_MEMORY

# CS0 Implementation
    implements CYGINT_HAL_KINETIS_FB_CS0
    implements CYGINT_DEVS_RAM0_MICRON_CELLULAR
    requires { is_active(CYGPKG_HAL_CORTEXM_KINETIS_FBRAM) implies
                         CYGHWR_HAL_KINETIS_FBR_SIZE == CYGHWR_HAL_KINETIS_FB_CS0_SIZE }

    cdl_option CYGHWR_HAL_KINETIS_FB_CS0_AR {
        display "Base address"
        flavor data
        parent CYGHWR_HAL_KINETIS_FB_CS0
        default_value  0x60000000
    }

    cdl_option CYGHWR_HAL_KINETIS_FB_CS0_SIZE {
        display "Size \[Bytes\]"
        flavor data
        legal_values  { 0x00040000  0x00400000 CYGHWR_RAM0_MICRON_CELLULAR_SIZE }
        parent        CYGHWR_HAL_KINETIS_FB_CS0
        default_value CYGHWR_RAM0_MICRON_CELLULAR_SIZE
    }

    cdl_option CYGHWR_HAL_KINETIS_FB_CS0_BASE {
        display "Memory base address"
        flavor data
        parent CYGHWR_HAL_KINETIS_FB_CS0
        calculated CYGHWR_HAL_KINETIS_FB_CS0_AR
    }

    cdl_component CYGHWR_HAL_KINETIS_FB_CS0_MR {
        display "Mask register"
        flavor data
        parent CYGHWR_HAL_KINETIS_FB_CS0
        default_value 0x00FF0001

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_MR_WP {
            display "Write protect"
            flavor bool
            default_value 0
        }
    }

    cdl_component CYGHWR_HAL_KINETIS_FB_CS0_CR {
        display "Control register"
        flavor none
        parent CYGHWR_HAL_KINETIS_FB_CS0

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_WS {
            display "Wait states"
            flavor data
            default_value 3
            legal_values 0 to 63
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_BLS {
            display "Byte lane shift"
            flavor data
            legal_values { 0 1 }
            default_value 1
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_AA {
            display "Auto acknowledge enable"
            flavor data
            legal_values { 0 1 }
            default_value 1
        }

        cdl_component CYGHWR_HAL_KINETIS_FB_CS0_CR_PSB {
            display "Port size (bits)"
            flavor data
            legal_values { 32 8 16 "-16" }
            default_value 16

        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_SWSEN {
            display "Secondary wait states enable"
            flavor data
            legal_values { 0 1 }
            default_value 1
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_SWS {
            display "Secondary wait states"
            flavor data
            legal_values 0 to 63
            default_value 0

        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_EXALE {
            display "Extended address latch enable"
            flavor data
            legal_values { 0 1 }
            default_value 1
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_ASET {
            display "Address setup"
            flavor data
            legal_values { 0 1 2 3 }
            default_value 0
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_RDAH {
            display "Read address hold or deselect"
            flavor data
            legal_values { 0 1 2 3 }
            default_value 0
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_WRAH {
            display "Write address hold or deselect"
            flavor data
            legal_values { 0 1 2 3 }
            default_value 0
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_BEM {
            display "Byte enable mode"
            flavor data
            legal_values { 0 1 }
            default_value 1
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_BSTR {
            display "Burst read enable"
            flavor data
            legal_values { 0 1 }
            default_value 1
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_BSTW {
            display "Burst write enable"
            flavor data
            legal_values { 0 1 }
            default_value 0
        }
    }

    cdl_component CYGHWR_HAL_KINETIS_FB_CS0_CR_IS {
        display "Control register initial setting."
        flavor none
        parent CYGHWR_HAL_KINETIS_FB_CS0

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_IS_WS {
            display "Wait states"
            flavor data
            default_value 3
            legal_values 0 to 63
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_IS_AA {
            display "Auto acknowledge enable"
            flavor data
            legal_values { 0 1 }
            default_value 1
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_IS_SWSEN {
            display "Secondary wait states enable"
            flavor data
            legal_values { 0 1 }
            default_value 0
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_IS_SWS {
            display "Secondary wait states"
            flavor data
            legal_values 0 to 63
            default_value 0

        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_IS_EXALE {
            display "Extended address latch enable"
            flavor data
            legal_values { 0 1 }
            default_value 1
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_IS_ASET {
            display "Address setup"
            flavor data
            legal_values { 0 1 2 3 }
            default_value 0
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_IS_RDAH {
            display "Read address hold or deselect"
            flavor data
            legal_values { 0 1 2 3 }
            default_value 0
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_IS_WRAH {
            display "Write address hold or deselect"
            flavor data
            legal_values { 0 1 2 3 }
            default_value 0
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_IS_BEM {
            display "Byte enable mode"
            flavor data
            legal_values { 0 1 }
            default_value 1
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_IS_BSTR {
            display "Burst read enable"
            flavor data
            legal_values { 0 1 }
            default_value 0
        }

        cdl_option CYGHWR_HAL_KINETIS_FB_CS0_CR_IS_BSTW {
            display "Burst write enable"
            flavor data
            legal_values { 0 1 }
            default_value 0
        }
    }
# CS0 Implementation End
# FlexBus  Implementation End

    cdl_option CYGHWR_HAL_KINETIS_FB_EXTRAM_SIZE {
        display "External RAM size"
        flavor data
        calculated CYGHWR_HAL_KINETIS_FB_CS0_SIZE
    }

    cdl_option CYGHWR_HAL_KINETIS_FB_EXTRAM_BASE {
        display "External RAM base address"
        flavor data
        calculated CYGHWR_HAL_KINETIS_FB_CS0_BASE
    }

    cdl_option CYGHWR_FREESCALE_ENET_MII_MDC_HAL_CLOCK {
        display "ENET MII MDC clock provided by HAL"
        flavor data
        active_if CYGPKG_DEVS_ETH_FREESCALE_ENET
        parent CYGPKG_DEVS_ETH_FREESCALE_ENET
        calculated CYGHWR_HAL_CORTEXM_KINETIS_CLK_PER_BUS
        description "
            ENET needs a clock with typical frequency of up to 2.5 MHz for
            MII MDC. The input clock, typically provided by HAL, is further
            divided by ENET according to setting of ENET MSCR register in order to
            provide frequency within 2.5 MHz range."
     }

    cdl_option CYGHWR_HAL_FREESCALE_ENET_E0_1588_PORT {
        display "IEEE 1588 Port"
        active_if CYGSEM_DEVS_ETH_FREESCALE_ENET_1588
        parent CYGSEM_DEVS_ETH_FREESCALE_ENET_1588
        flavor data
        default_value { "B" }
        legal_values { "B" "C" "User" }
        description "
            Digital I/O provided by HAL for ENET IEEE 1588 timers."
    }



    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
        Global build options including control over
        compiler flags, linker flags and choice of toolchain."

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-eabi" }
            description "
            This option specifies the command prefix used when
            invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGBLD_GLOBAL_WARNFLAGS . "-mcpu=cortex-m3 -mthumb -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions" }
            description   "
            This option controls the global compiler flags which are used to
            compile all packages by default. Individual packages may define
            options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-mcpu=cortex-m3 -mthumb -Wl,--gc-sections -Wl,-static -Wl,-n -g -nostdlib" }
            description   "
            This option controls the global linker flags. Individual
            packages may define options which override these global flags."
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        requires      { CYGDBG_HAL_CRCTABLE_LOCATION == "ROM" }
        description   "
        Enable this option if this program is to be used as a ROM monitor,
        i.e. applications will be loaded into RAM on the board, and this
        ROM monitor may process exceptions or interrupts generated from the
        application. This enables features such as utilizing a separate
        interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
        display       "Work with a ROM monitor"
        flavor        booldata
        legal_values  { "Generic" "GDB_stubs" }
        default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "RAM" }
        description   "
        Support can be enabled for different varieties of ROM monitor.
        This support changes various eCos semantics such as the encoding
        of diagnostic output, or the overriding of hardware interrupt
        vectors.
        Firstly there is \"Generic\" support which prevents the HAL
        from overriding the hardware vectors that it does not use, to
        instead allow an installed ROM monitor to handle them. This is
        the most basic support which is likely to be common to most
        implementations of ROM monitor.
        \"GDB_stubs\" provides support when GDB stubs are included in
        the ROM monitor or boot ROM."
    }

    cdl_component CYGBLD_HAL_CORTEXM_TWR_MK60N512_GDB_STUBS {
        display "Create StubROM SREC and binary files"
        active_if CYGBLD_BUILD_COMMON_GDB_STUBS
        no_define
        calculated 1
        requires { CYG_HAL_STARTUP == "ROM" }

        make -priority 325 {
            <PREFIX>/bin/stubrom.srec : <PREFIX>/bin/gdb_module.img
            $(OBJCOPY) -O srec $< $@
        }
        make -priority 325 {
            <PREFIX>/bin/stubrom.bin : <PREFIX>/bin/gdb_module.img
            $(OBJCOPY) -O binary $< $@
        }

        description "This component causes the ELF image generated by the
        build process to be converted to S-Record and binary
        files."
    }
}
