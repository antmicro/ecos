
# ====================================================================
#
#      hal_arm_mac7100_mace1.cdl
#
#      ARM MAC7100 MACE1 HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003, 2006 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Ilija Koco <ilijak@siva.com.mk>
# Contributors:   
# Date:           2006-04-12
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_MAC7100_MACE1 {
    display       "MACE1 - MAC7100 eval board HAL"
    parent        CYGPKG_HAL_ARM_MAC7100
    define_header hal_arm_mac7100_mace1.h
    include_dir   cyg/hal
    hardware
    description   "
        The MACE1 HAL package provides the support needed to run
        eCos on an MACE1 - MAC7100 eval board."

    compile       mace1_misc.c

    requires      { CYGHWR_HAL_ARM_MAC7100 == "MAC7121" }
    requires      { CYGNUM_PIT_CHAN_CLOCK_PRIORITY == 
                    CYGNUM_KERNEL_COUNTERS_CLOCK_ISR_PRIORITY }

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_arm_mac7100.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_mac7100_mace1.h>"
        puts $::cdl_header "#define HAL_PLATFORM_CPU    \"ARM7TDMI\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Freescale MAC7100/MACE1\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
    }

    cdl_component CYG_PIT_CLOCKS {
        display "Real time clock configuration."
        flavor   none
        description "
            Periodic Interrupt Timer Module - PIT comprizes 11 timer
            channels.  RTI channel (PIT0) as well as PIT1 .. PIT4 can
            generate interrupts and are eligible for the real time
            clock.  "

        cdl_option CYGNUM_PIT_CHAN_CLOCK {
            display      "System CLOCK device"
            flavor       data
            legal_values 0 to 4
            default_value   3
            requires {CYGNUM_PIT_CHAN_CLOCK != CYGNUM_PIT_CHAN_US}
            description "
                RTI (PIT0) and PIT1 .. PIT4 can be used for ral time
                clock.  RTI is clocked by oscillator clock while
                channels 1 to 4 by 1/2 system clock frequency.
                Selection of RTI vs PIT1 .. PIT4 affects Real-time
                clock period (see Real-time clock constants).  NOTE:
                Real time clock channel must not be the same as US
                delay channel.
            "
        }

        cdl_option CYGNUM_PIT_CHAN_CLOCK_PRIORITY {
            display      "System clock's INTC priority"
            flavor       data
            legal_values 0 to 15
            default_value   12
            description "
                INTC has 16 interrupt levels: 0 (lowest) to 15 (highest).
            "
        }

        cdl_option CYGNUM_PIT_CHAN_US {
            display      "PIT channel for us delay"
            flavor       data
            legal_values 0 to 4
            default_value   0
            requires {CYGNUM_PIT_CHAN_CLOCK != CYGNUM_PIT_CHAN_US}
            description "
                RTI is clocked by oscillator while channels PIT1
                .. PIT4 by half system clock frequency, hence RTI
                should allow for larger maximal period.  NOTE: US
                delay channel must not be the same as real time clock
                channel.
            "
        }
    }
    
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none

        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            default_value 1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            default_value (CYGNUM_PIT_CHAN_CLOCK !=0 ? \
                (CYGNUM_HAL_ARM_MAC7100_CLOCK_SPEED / 2 / CYGNUM_HAL_RTC_DENOMINATOR - 1) : \
                (CYGNUM_HAL_ARM_MAC7100_Q_FREQ / CYGNUM_HAL_RTC_DENOMINATOR - 1))
        }
    }
    
    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        calculated {"ROM"}
        no_define
        define -file system.h CYG_HAL_STARTUP
        description   "
            Current MACE1 port supports only ROM startup type."
    }

    # Real-time clock/counter specifics

    cdl_component CYG_HAL_MAC7100_OSC {
        display "System Clocks Module"
        flavor  none

        cdl_option CYGNUM_HAL_ARM_MAC7100_F_OSC {
            display       "FOSC - Oscillator clock"
            flavor        data
            default_value 8000000
        }
        
        cdl_option CYGNUM_HAL_ARM_MAC7100_FDIV {
            display       "FDIV - Frequency divider for PLL"
            flavor        booldata
            legal_values 0 to 16
            default_value 2
            description "
                If enabled (FDIV != 0), 
                   you set divider for PLL. 
                   Then REFDV is calculated as REFDV=FDIV-1;
                If disabled (FDIV == 0), 
                   REFDV is calculated from FOSC so that referent frequency 
                   for PLL is 500kHz.
                   SYNR is then derived from desired CPU clock, FOSC and REFDV.
                "
        }
    }

    cdl_option CYGNUM_HAL_ARM_MAC7100_CLOCK_SPEED {
        display       "CPU clock - PLL frequency"
        flavor        data
        default_value 48000000
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        legal_values 0 1 2
        default_value   2
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The MAC7100 MACE1 board has two serial ports. This option
            chooses which port will be used to connect to a host
            running GDB."
     }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    0
         description      "
            The MAC7100 MACE1 board has two serial ports. This option
            chooses which port will be used for diagnostic output."
     }
     
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400
        default_value 38400
        description   "
            This option selects the baud rate used for the diagnostic port."
    }
 
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
         display       "GDB serial port baud rate"
         flavor        data
         legal_values  9600 19200 38400
         default_value 38400
         description   "
            This option controls the baud rate used for the GDB connection."
     }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" || 
                        CYG_HAL_STARTUP == "ROMRAM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "Generic" "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             Firstly there is \"Generic\" support which prevents the HAL
             from overriding the hardware vectors that it does not use, to
             instead allow an installed ROM monitor to handle them. This is
             the most basic support which is likely to be common to most
             implementations of ROM monitor.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
     }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to a binary image suitable for ROM programming."
    
            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }

        }
    }
 
    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
        Global build options including control over
        compiler flags, linker flags and choice of toolchain."

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-eabi"}
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGBLD_GLOBAL_WARNFLAGS . CYGBLD_ARCH_CFLAGS .
                            "-mcpu=arm7tdmi -gdwarf-2 -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions " }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define options which
                override these global flags."

        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { CYGBLD_ARCH_LDFLAGS . "-mcpu=arm7tdmi -Wl,--gc-sections -Wl,-static -gdwarf-2 -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { (CYG_HAL_STARTUP == "RAM") ?    "arm_mac7100_mace1_ram" :
                     (CYG_HAL_STARTUP == "ROMRAM") ? "arm_mac7100_mace1_romram" :
                                                     "arm_mac7100_mace1_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { (CYG_HAL_STARTUP == "RAM") ? "<pkgconf/mlt_arm_mac7100_mace1_ram.ldi>" :
                         (CYG_HAL_STARTUP == "ROMRAM") ? "<pkgconf/mlt_arm_mac7100_mace1_romram.ldi>" :
                                                      "<pkgconf/mlt_arm_mac7100_mace1_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { (CYG_HAL_STARTUP == "RAM") ? "<pkgconf/mlt_arm_mac7100_mace1_ram.h>" :
                         (CYG_HAL_STARTUP == "ROMRAM") ? "<pkgconf/mlt_arm_mac7100_mace1_romram.h>" :
                                                      "<pkgconf/mlt_arm_mac7100_mace1_rom.h>" }
        }
    }
}
