# ====================================================================
#
#      hal_sh_sh3.cdl
#
#      SH3 variant HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  jskov
# Contributors:
# Date:           2000-10-30
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_SH_SH3 {
    display       "SH3 variant"
    parent        CYGPKG_HAL_SH
    hardware
    include_dir   cyg/hal
    define_header hal_sh_sh3.h
    description   "
        The SH3 (SuperH 3) variant HAL package provides generic
        support for SH3 variant CPUs."

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H   <pkgconf/hal_sh_sh3.h>"
        puts $::cdl_header "#define CYGBLD_HAL_VAR_EXCEPTION_MODEL_H   <cyg/hal/hal_var_bank.h>"
        puts $::cdl_header "#define CYGBLD_HAL_VAR_EXCEPTION_MODEL_INC <cyg/hal/hal_var_bank.inc>"
        puts $::cdl_header "#define CYGBLD_HAL_VAR_INTR_MODEL_H   <cyg/hal/hal_intr_excevt.h>"
    }

    compile       sh3_sci.c sh3_scif.c var_misc.c variant.S

    # The "-o file" is a workaround for CR100958 - without it the
    # output file would end up in the source directory under CygWin.
    # n.b. grep does not behave itself under win32
    make -priority 1 {
        <PREFIX>/include/cyg/hal/sh3_offsets.inc : <PACKAGE>/src/var_mk_defs.c
        $(CC) $(ACTUAL_CFLAGS) $(INCLUDE_PATH) -Wp,-MD,sh3_offsets.tmp -o var_mk_defs.tmp -S $<
        fgrep .equ var_mk_defs.tmp | sed s/#// > $@
        @echo $@ ": \\" > $(notdir $@).deps
        @tail -n +2 sh3_offsets.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm sh3_offsets.tmp var_mk_defs.tmp
    }

    # CPU variant supported
    cdl_option CYGPKG_HAL_SH_7707A {
        display       "SH 7707A microprocessor"
        parent        CYGPKG_HAL_SH_CPU
        implements    CYGINT_HAL_SH_VARIANT
        implements    CYGINT_HAL_SH_CPG_T2
        default_value 0
        no_define
        define        -file=system.h CYGPKG_HAL_SH_7707A
        description "
            The SH3 7707A microprocessor. This is an embedded part that in
            addition to the SH3 processor core has built in peripherals
            such as memory controllers, serial ports, LCD controller and
            timers/counters."               
        define_proc {
            puts $cdl_system_header "#define CYGBLD_HAL_CPU_MODULES_H <cyg/hal/mod_7707a.h>"
        }
    }
    
    cdl_option CYGPKG_HAL_SH_7708 {
        display       "SH 7708 microprocessor"
        parent        CYGPKG_HAL_SH_CPU
        implements    CYGINT_HAL_SH_VARIANT
        implements    CYGINT_HAL_SH_CPG_T1
        default_value 0
        no_define
        define        -file=system.h CYGPKG_HAL_SH_7708
        description "
            The SH3 7708 microprocessor. This is an embedded part that in
            addition to the SH3 processor core has built in peripherals
            such as memory controllers, serial ports and
            timers/counters."               
        define_proc {
            puts $cdl_system_header "#define CYGBLD_HAL_CPU_MODULES_H <cyg/hal/mod_7708.h>"
        }
    }
    
    cdl_option CYGPKG_HAL_SH_7709A {
        display       "SH 7709A microprocessor"
        parent        CYGPKG_HAL_SH_CPU
        implements    CYGINT_HAL_SH_VARIANT
        implements    CYGINT_HAL_SH_CPG_T3
        implements    CYGINT_HAL_SH_DMA_CHANNELS
        implements    CYGINT_HAL_SH_DMA_CHANNELS
        implements    CYGINT_HAL_SH_DMA_CHANNELS
        implements    CYGINT_HAL_SH_DMA_CHANNELS
        default_value 1
        no_define
        define        -file=system.h CYGPKG_HAL_SH_7709A
        description "
            The SH3 7709A microprocessor. This is an embedded part that in
            addition to the SH3 processor core has built in peripherals
            such as memory controllers, DMA controllers, A/D and D/A
            converters, serial ports and timers/counters."               
        define_proc {
            puts $cdl_system_header "#define CYGBLD_HAL_CPU_MODULES_H <cyg/hal/mod_7709a.h>"
        }
    }

    cdl_option CYGPKG_HAL_SH_7709R {
        display       "SH 7709R microprocessor"
        parent        CYGPKG_HAL_SH_CPU
        implements    CYGINT_HAL_SH_VARIANT
        implements    CYGINT_HAL_SH_CPG_T3
        default_value 0
        no_define
        define        -file=system.h CYGPKG_HAL_SH_7709R
        description "
            The SH3 7709R microprocessor. This is an embedded part that in
            addition to the SH3 processor core has built in peripherals
            such as memory controllers, DMA controllers, A/D and D/A
            converters, serial ports and timers/counters."               
        define_proc {
            puts $cdl_system_header "#define CYGBLD_HAL_CPU_MODULES_H <cyg/hal/mod_7709r.h>"
        }
    }

    cdl_option CYGPKG_HAL_SH_7709S {
        display       "SH 7709S microprocessor"
        parent        CYGPKG_HAL_SH_CPU
        implements    CYGINT_HAL_SH_VARIANT
        implements    CYGINT_HAL_SH_CPG_T3
        implements    CYGINT_HAL_SH_DMA_CHANNELS
        implements    CYGINT_HAL_SH_DMA_CHANNELS
        implements    CYGINT_HAL_SH_DMA_CHANNELS
        implements    CYGINT_HAL_SH_DMA_CHANNELS
        default_value 0
        no_define
        define        -file=system.h CYGPKG_HAL_SH_7709S
        description "
            The SH3 7709S microprocessor. This is an embedded part that in
            addition to the SH3 processor core has built in peripherals
            such as memory controllers, DMA controllers, A/D and D/A
            converters, serial ports and timers/counters."               
        define_proc {
            puts $cdl_system_header "#define CYGBLD_HAL_CPU_MODULES_H <cyg/hal/mod_7709s.h>"
        }
    }
    
    cdl_option CYGPKG_HAL_SH_7729 {
        display       "SH 7729 microprocessor"
        parent        CYGPKG_HAL_SH_CPU
        implements    CYGINT_HAL_SH_VARIANT
        implements    CYGINT_HAL_SH_CPG_T3
        default_value 0
        no_define
        define        -file=system.h CYGPKG_HAL_SH_7729
        description "
            The SH3 7729 microprocessor. This is an embedded part that in
            addition to the SH3 processor core has built in peripherals
            such as memory controllers, serial ports, and timers/counters,
            and a DSP engine."
        define_proc {
            puts $cdl_system_header "#define CYGBLD_HAL_CPU_MODULES_H <cyg/hal/mod_7729.h>"
        }
    }
    
    cdl_component CYGHWR_HAL_SH_CLOCK_SETTINGS {
        display          "SH on-chip generic clock controls"
        description      "
            The various clocks used by the system are controlled by
            these options, some of which are derived from platform
            settings."
        flavor        none
        no_define

        cdl_interface CYGINT_HAL_SH_CPG_T1 {
            display     "Clock pulse generator type 1"
        }

        cdl_interface CYGINT_HAL_SH_CPG_T2 {
            display     "Clock pulse generator type 2"
        }

        cdl_interface CYGINT_HAL_SH_CPG_T3 {
            display     "Clock pulse generator type 3"
        }


        cdl_option CYGHWR_HAL_SH_TMU_PRESCALE_0 {
            display       "TMU counter 0 prescaling"
            description   "
                The peripheral clock is driving the counter used for
                the real-time clock, prescaled by this factor."
            flavor        data
            legal_values  { 4 16 64 256 }
            default_value 4
        }

        cdl_option CYGHWR_HAL_SH_RTC_PRESCALE {
            display       "eCos RTC prescaling"
            flavor        data
            calculated    CYGHWR_HAL_SH_TMU_PRESCALE_0
        }

        cdl_option CYGHWR_HAL_SH_CLOCK_CKIO {
            display    "CKIO clock"
            no_define
            flavor     data
            # CKIO is either XTAL or PLL2 output
            calculated { CYGINT_HAL_SH_CPG_T1 ? (
                             (CYGHWR_HAL_SH_OOC_CLOCK_MODE == 7) 
                             ? (CYGHWR_HAL_SH_OOC_XTAL)
                             : CYGHWR_HAL_SH_PLL2_OUTPUT
                         )
                         : CYGINT_HAL_SH_CPG_T2 ? (
                             (CYGHWR_HAL_SH_OOC_CLOCK_MODE == 2) 
                             ? (CYGHWR_HAL_SH_OOC_XTAL)
                             : CYGHWR_HAL_SH_PLL2_OUTPUT
                         )
                         : CYGINT_HAL_SH_CPG_T3 ? (
                             (CYGHWR_HAL_SH_OOC_CLOCK_MODE == 7) 
                             ? (CYGHWR_HAL_SH_OOC_XTAL)
                             : CYGHWR_HAL_SH_PLL2_OUTPUT
                         )
                         : 0 }
        }

        cdl_option CYGHWR_HAL_SH_PLL1_OUTPUT {
            display    "The clock output from PLL1"
            no_define
            flavor     data
            calculated { CYGHWR_HAL_SH_CLOCK_CKIO * CYGHWR_HAL_SH_OOC_PLL_1 }
        }

        cdl_option CYGHWR_HAL_SH_PLL2_OUTPUT {
            display    "The clock output from PLL2"
            no_define
            flavor     data
            calculated { CYGINT_HAL_SH_CPG_T1 ? (
                             (CYGHWR_HAL_SH_OOC_XTAL * CYGHWR_HAL_SH_OOC_PLL_2)
                         )
                         : CYGINT_HAL_SH_CPG_T2 ? (
                             (CYGHWR_HAL_SH_OOC_CLOCK_MODE == 5)
                             ? (CYGHWR_HAL_SH_OOC_XTAL / 2)
                             : (CYGHWR_HAL_SH_OOC_CLOCK_MODE == 6) 
                             ? (14745600)
                             : (CYGHWR_HAL_SH_OOC_CLOCK_MODE == 7) 
                             ? (11075600)
                             : (CYGHWR_HAL_SH_OOC_XTAL * CYGHWR_HAL_SH_OOC_PLL_2)
                         )
                         : CYGINT_HAL_SH_CPG_T3 ? (
                             (CYGHWR_HAL_SH_OOC_XTAL * CYGHWR_HAL_SH_OOC_PLL_2)
                         )
                         : 0 }
        }


        cdl_option CYGHWR_HAL_SH_DIVIDER1_INPUT {
            display    "The clock input to divider 1"
            no_define
            flavor     data
            # DIV1 input is either PLL2 output or PLL1 output
            calculated { (CYGHWR_HAL_SH_OOC_PLL_1 == 0)
                           ? CYGHWR_HAL_SH_PLL2_OUTPUT
                           : CYGHWR_HAL_SH_PLL1_OUTPUT }
        }

        cdl_option CYGHWR_HAL_SH_DIVIDER2_INPUT {
            display    "The clock input to divider 2"
            no_define
            flavor     data
            # DIV2 input is either PLL2 output or PLL1 output
            calculated { CYGINT_HAL_SH_CPG_T1 ? (
                             (CYGHWR_HAL_SH_OOC_CLOCK_MODE == 3 || CYGHWR_HAL_SH_OOC_CLOCK_MODE == 4)
                             ? CYGHWR_HAL_SH_PLL2_OUTPUT
                             : CYGHWR_HAL_SH_PLL1_OUTPUT
                         )
                         : CYGINT_HAL_SH_CPG_T2 ? (
                             (CYGHWR_HAL_SH_OOC_CLOCK_MODE <= 2)
                             ? CYGHWR_HAL_SH_PLL1_OUTPUT
                             : CYGHWR_HAL_SH_PLL2_OUTPUT
                         )
                         : CYGINT_HAL_SH_CPG_T3 ? (
                             (CYGHWR_HAL_SH_OOC_CLOCK_MODE == 3 || CYGHWR_HAL_SH_OOC_CLOCK_MODE == 4)
                             ? CYGHWR_HAL_SH_PLL2_OUTPUT
                             : CYGHWR_HAL_SH_PLL1_OUTPUT
                         )
                         : 0 }
        }

        cdl_option CYGHWR_HAL_SH_PROCESSOR_SPEED {
            display          "Processor clock speed (MHz)"
            flavor           data
            calculated       { CYGHWR_HAL_SH_DIVIDER1_INPUT / CYGHWR_HAL_SH_OOC_DIVIDER_1 }
            description      "
                The core (CPU, cache and MMU) speed is computed from
                the input clock speed and the divider 1 setting."
        }

        cdl_option CYGHWR_HAL_SH_BOARD_SPEED {
            display          "Platform bus clock speed (MHz)"
            flavor           data
            calculated       { CYGHWR_HAL_SH_CLOCK_CKIO }
            description      "
                The platform bus speed is CKIO."
        }

        cdl_option CYGHWR_HAL_SH_ONCHIP_PERIPHERAL_SPEED {
            display          "Processor on-chip peripheral clock speed (MHz)"
            flavor           data
            calculated       { CYGHWR_HAL_SH_DIVIDER2_INPUT / CYGHWR_HAL_SH_OOC_DIVIDER_2 }
            description      "
                The peripheral speed is computed from the input clock
                speed and the divider 2 settings."
        }
    }

    cdl_option CYGNUM_HAL_SH_SH3_SCI_BAUD_RATE {
        display          "SCI serial port default baud rate"
        flavor data
        legal_values     { 4800 9600 14400 19200 38400 57600 115200 }
        default_value    { CYGNUM_HAL_SH_SH3_SCI_BAUD_RATE_DEFAULT ? \
                           CYGNUM_HAL_SH_SH3_SCI_BAUD_RATE_DEFAULT : 38400 }
        description      "
           This controls the default baud rate used for communicating
           with GDB / displaying diagnostic output."
    }

    cdl_option CYGNUM_HAL_SH_SH3_SCIF_BAUD_RATE {
        display          "SCIF serial ports default baud rate"
        flavor data
        legal_values     { 4800 9600 14400 19200 38400 57600 115200 }
        default_value    { CYGNUM_HAL_SH_SH3_SCIF_BAUD_RATE_DEFAULT ? \
                           CYGNUM_HAL_SH_SH3_SCIF_BAUD_RATE_DEFAULT : 38400 }
        description      "
           This controls the default baud rate used for communicating
           with GDB / displaying diagnostic output."
    }

    cdl_component CYGPKG_HAL_SH_INTERRUPT {
        display          "Interrupt controls"
        flavor     none
        no_define
        description      "
            Initial interrupt settings can be specified using these option."

        cdl_option CYGHWR_HAL_SH_IRQ_HANDLE_SPURIOUS_INTERRUPTS {
            display          "Handle spurious interrupts"
            default_value    0
            description      "
               The SH3 may generate spurious interrupts with INTEVT = 0
               when changing the BL bit of the status register. Enabling
               this option will cause such interrupts to be identified
               very early in the interrupt handler and be ignored.  Given
               that the SH HAL uses the I-mask to control interrupts,
               these spurious interrupts should not occur, and so there
               should be no reason to include the special handling code."
        }

        cdl_option CYGHWR_HAL_SH_IRQ_USE_IRQLVL {
            display          "Use IRQ0-3 pins as IRL input"
            default_value    0
            description      "
                It is possible for the IRQ0-3 pins to be used as IRL
                inputs by enabling this option."
        }

        cdl_option CYGHWR_HAL_SH_IRQ_ENABLE_IRLS_INTERRUPTS {
            display          "Enable IRLS interrupt pins"
            default_value    0
            active_if        CYGHWR_HAL_SH_IRQ_USE_IRQLVL
            description      "
                IRLS interrupt pins must be specifically
                activated. When they are, they will cause the same
                type of interrupt as those caused by the IRL pins. If
                IRL and IRLS pins signal an interrupt at the same
                time, the highest level interrupt will be generated.
                Only available on some cores, and probably share pins
                with other interrupt sources (PINT) which cannot be
                used in this configuration."
        }
    }

    # Cache settings
    cdl_option CYGHWR_HAL_SH_CACHE_MODE_P0 {
        display       "Select cache mode set for P0/U0/P3 at startup"
        parent        CYGPKG_HAL_SH_CACHE
        default_value { "WRITE_BACK" }
        legal_values  { "WRITE_BACK" "WRITE_THROUGH" }
        flavor        data
        description "
            Controls what cache mode the cache should be put in at
            startup for areas P0, U0 and P3. Write-back mode improves
            performance by letting dirty data to be kept in the
            cache for a period of time, allowing mutiple writes to
            the same cache line to be written back to memory in
            one memory transaction. In Write-through mode, each
            individual write will cause a memory transaction."
    }
    
    cdl_option CYGHWR_HAL_SH_CACHE_MODE_P1 {
        display       "Select cache mode set for P1 at startup"
        parent        CYGPKG_HAL_SH_CACHE
        default_value { "WRITE_BACK" }
        legal_values  { "WRITE_BACK" "WRITE_THROUGH" }
        flavor        data
        description "
            Controls what cache mode the cache should be put in at
            startup for area P1. Write-back mode improves
            performance by letting dirty data to be kept in the
            cache for a period of time, allowing mutiple writes to
            the same cache line to be written back to memory in
            one memory transaction. In Write-through mode, each
            individual write will cause a memory transaction."
    }
}
