# ====================================================================
#
#      fec_eth_drivers.cdl
#
#      Ethernet drivers - platform dependent support for PowerPC MPC8260
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      mtek
# Original data:  gthomas
# Contributors:
# Date:           2002-02-20
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_POWERPC_QUICC2 {
    display       "MPC8260 FEC ethernet driver"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_HAL_POWERPC 
    active_if	  CYGPKG_HAL_POWERPC_MPC8260

    implements    CYGHWR_NET_DRIVERS
    implements    CYGHWR_NET_DRIVER_ETH0
    include_dir   .
    include_files ; # none _exported_ whatsoever

    description   "Fast ethernet driver for PowerPC MPC8260 boards."
    compile       -library=libextras.a if_fec.c EnetPHY.c

    cdl_option CYGNUM_DEVS_ETH_POWERPC_QUICC2_BUFSIZE {
        display       "Buffer size"
        flavor        data
        default_value 1540
        description   "
            This option specifies the size of the internal buffers used
            for the PowerPC FEC/ethernet device."
    }

    cdl_option CYGNUM_DEVS_ETH_POWERPC_QUICC2_TxNUM {
        display       "Number of output buffers"
        flavor        data
        legal_values  2 to 16
        default_value 4
        description   "
            This option specifies the number of output buffer packets
            to be used for the PowerPC FEC/ethernet device."
    }

    cdl_option CYGNUM_DEVS_ETH_POWERPC_QUICC2_RxNUM {
        display       "Number of input buffers"
        flavor        data
        legal_values  2 to 16
        default_value 4
        description   "
            This option specifies the number of input buffer packets
            to be used for the PowerPC FEC/ethernet device."
    }

    cdl_component CYGPKG_DEVS_ETH_POWERPC_QUICC2_OPTIONS {
        display "MPC8260 FEC ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_POWERPC_QUICC2_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the MPC8260 FEC ethernet driver package. 
		These flags are used in addition to the set of global 
		flags."
        }
    }
}
