# ====================================================================
#
#      i386_pc_rltk8139_eth_drivers.cdl
#
#      Ethernet drivers - support for RealTek 8139 ethernet controller
#      on i386 PC target
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Eric Doenges
# Contributors:
# Date:           2003-07-16
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_I386_PC_RLTK8139 {
    display       "PC RealTek 8139 ethernet driver"
    description   "Ethernet driver for standard PC's."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_HAL_I386_PC

    include_dir   cyg/io

    # FIXME: This really belongs in the RealTek_8139 package ?
    cdl_interface CYGINT_DEVS_ETH_RLTK_8139_REQUIRED {
        display   "RealTek 8139 ethernet driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_RLTK_8139_INL <cyg/io/devs_eth_i386_pc_rltk8139.inl>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_RLTK_8139_CFG <pkgconf/devs_eth_i386_pc_rltk8139.h>"
        puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
    }

    cdl_component CYGPKG_DEVS_ETH_I386_PC_RLTK8139_ETH0 {
        display       "Ethernet port 0 driver"
        flavor        bool
        default_value 1

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH0
        implements CYGINT_DEVS_ETH_RLTK_8139_REQUIRED

        cdl_option CYGDAT_DEVS_ETH_I386_PC_RLTK8139_ETH0_NAME {
            display       "Device name for the ETH0 ethernet port 0 driver"
            flavor        data
            default_value {"\"eth0\""}
            description   "
                This option sets the name of the ethernet device for the
                RealTek 8139 ethernet port 0."
        }
    }

    cdl_component CYGPKG_DEVS_ETH_I386_PC_RLTK8139_ETH1 {
        display       "Ethernet port 1 driver"
        flavor        bool
        default_value 0

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH1
        implements CYGINT_DEVS_ETH_RLTK_8139_REQUIRED

        cdl_option CYGDAT_DEVS_ETH_I386_PC_RLTK8139_ETH1_NAME {
            display       "Device name for the ETH1 ethernet port 1 driver"
            flavor        data
            default_value {"\"eth1\""}
            description   "
                This option sets the name of the ethernet device for the
                RealTek 8139 ethernet port 1."
        }
    }
}
