##==========================================================================
##
##      hal_cortexm_stm32.cdl
##
##      Cortex-M STM32 variant HAL configuration data
##
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008, 2011 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##==========================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):    nickg
## Contributors: jld
## Date:         2008-07-30
##
######DESCRIPTIONEND####
##
##==========================================================================

cdl_package CYGPKG_HAL_CORTEXM_STM32 {
    display       "Cortex-M3/-M4/-M7 STM32 Variant"
    parent        CYGPKG_HAL_CORTEXM
    hardware
    include_dir   cyg/hal
    define_header hal_cortexm_stm32.h
    description   "
        This package provides generic support for the ST Cortex-M based STM32
        microcontroller family.
        It is also necessary to select a variant and platform HAL package."

    compile       hal_diag.c stm32_misc.c stm32_dma.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_VIRTUAL_VECTOR_COMM_BAUD_SUPPORT
    implements    CYGINT_PROFILE_HAL_TIMER

    requires      { (CYGHWR_HAL_CORTEXM == "M3") || (CYGHWR_HAL_CORTEXM == "M4") || (CYGHWR_HAL_CORTEXM == "M7") }

    cdl_component CYGHWR_HAL_CORTEXM_STM32_SELECTION {
        display          "STM32 processor selection"
        no_define
        flavor           none
        description      "
            The options within this component allow you to select which STM32
            processor is in use."


    cdl_option CYGHWR_HAL_CORTEXM_STM32 {
            display          "STM32 processor variant in use"
        flavor           data
            default_value    { (CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F1") ? CYGHWR_HAL_CORTEXM_STM32_F1 : \
                               (CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F2") ? CYGHWR_HAL_CORTEXM_STM32_F2 : \
                               (CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F7") ? CYGHWR_HAL_CORTEXM_STM32_F7 : \
			       CYGHWR_HAL_CORTEXM_STM32_F4 }
            # At some point we'll add the L1, etc. here.
        description      "The STM32 has several variants, the main differences
                          being in the size of on-chip FLASH and SRAM
                          and numbers of some peripherals. This option
                          allows the platform HAL to select the specific
                          microcontroller fitted."
    }

        cdl_option CYGHWR_HAL_CORTEXM_STM32_FAMILY {
            display          "Processor family in use"
            flavor           data
            default_value    { "F1" }
            legal_values     { "F1" "F2" "F4" "F7" }
	    # NOTE: F1/F2 imply CYGHWR_HAL_CORTEXM_M3 and F4 implies CYGHWR_HAL_CORTEXM_M4
            description      "
                Which family of STM32 processors is in use. This will
                usually be the leading part of the processor model name."
        }

	# NOTE: This allows later L1 support to still select "FAMILY_HIPERFORMANCE" if the I/O is the same:
        cdl_option CYGHWR_HAL_CORTEXM_STM32_FAMILY_HIPERFORMANCE {
            display     "Part belongs to ST Hi-Performance family"
	    active_if   { (CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F2") || (CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F4" || CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F7") }
	    calculated  { (CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F2") || (CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F4" || CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F7") }
            description "
	        Indicates that this part conforms to the I/O
		definitions for the Hi-Performance family of
		devices. Currently this includes the STM32 F2 and F4
		devices."
        }

        cdl_option CYGHWR_HAL_CORTEXM_STM32_F1 {
            display          "F1 processor family selection"
            flavor           data
            active_if        { CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F1" }
            default_value    {"F103ZE"}
            legal_values     {"F103RC" "F103VC" "F103ZC"
                              "F103RD" "F103VD" "F103ZD"
                              "F103RE" "F103VE" "F103ZE"
                              "F105R8" "F105V8"
                              "F105RB" "F105VB"
                              "F105RC" "F105VC"
                              "F107RB" "F107VB"
                              "F107RC" "F107VC"
                             }
            requires         { CYGHWR_HAL_CORTEXM_STM32 == CYGHWR_HAL_CORTEXM_STM32_F1 }
            description "
                This option specifies which member of the STM32F1 family is
                in use."
        }

        cdl_option CYGHWR_HAL_CORTEXM_STM32_F2 {
            display          "F2 processor family selection"
            flavor           data
            active_if        { CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F2" }
            default_value    {"F207IG"}
            legal_values     {"F205RB" "F205RC" "F205RE" "F205RF" "F205RG"
                              "F205VB" "F205VC" "F205VE" "F205VF" "F205VG"
                              "F205ZB" "F205ZC" "F205ZE" "F205ZF" "F205ZG"
                              "F207VB" "F207VC" "F207VE" "F207VF" "F207VG"
                              "F207ZB" "F207ZC" "F207ZE" "F207ZF" "F207ZG"
                              "F207IB" "F207IC" "F207IE" "F207IF" "F207IG"
                             }
            requires         { CYGHWR_HAL_CORTEXM_STM32 == CYGHWR_HAL_CORTEXM_STM32_F2 }
            description "
                This option specifies which member of the STM32F2 family is
                in use."
        }

        cdl_option CYGHWR_HAL_CORTEXM_STM32_F4 {
            display          "F4 processor family selection"
            flavor           data
            active_if        { CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F4" }
            default_value    {"F407IG"}
            # NOTEs: The "F4xxxE" parts have 512MB on-chip flash and
            # the "F4xxxG" parts have 1MB on-chip flash. The "F41xxx"
            # parts have CRYPTO support.
            legal_values     {"F405RG" "F405VG" "F405ZG"
                              "F415RG" "F415VG" "F415ZG"
                              "F407IG" "F407VG" "F407ZG"
                              "F407IE" "F407VE" "F407ZE"
                              "F417IG" "F417VG" "F417ZG"
                              "F417IE" "F417VE" "F417ZE"
                             }
            requires         { CYGHWR_HAL_CORTEXM_STM32 == CYGHWR_HAL_CORTEXM_STM32_F4 }
            description "
                This option specifies which member of the STM32F4 family is
                in use."
        }

        cdl_option CYGHWR_HAL_CORTEXM_STM32_F7 {
            display          "F7 processor family selection"
            flavor           data
            active_if        { CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F7" }
            default_value    {"F707IG"}
	    # NOTES: Copy from STM32_F4
            legal_values     {"F705RG" "F705VG" "F705ZG"
                              "F715RG" "F715VG" "F715ZG"
                              "F707IG" "F707VG" "F707ZG"
                              "F707IE" "F707VE" "F707ZE"
                              "F717IG" "F717VG" "F717ZG"
                              "F717IE" "F717VE" "F717ZE"
                             }
            requires         { CYGHWR_HAL_CORTEXM_STM32 == CYGHWR_HAL_CORTEXM_STM32_F7 }
            description "
                This option specifies which member of the STM32F7 family is
                in use."
        }
    }

    cdl_option CYGHWR_HAL_CORTEXM_STM32_CONNECTIVITY {
        display         "Part belongs to connectivity family"
        default_value   { (CYGHWR_HAL_CORTEXM_STM32 == "F105R8") || (CYGHWR_HAL_CORTEXM_STM32 == "F105V8") ||
                          (CYGHWR_HAL_CORTEXM_STM32 == "F105RB") || (CYGHWR_HAL_CORTEXM_STM32 == "F105VB") ||
                          (CYGHWR_HAL_CORTEXM_STM32 == "F105RC") || (CYGHWR_HAL_CORTEXM_STM32 == "F105VC") ||
                          (CYGHWR_HAL_CORTEXM_STM32 == "F107RB") || (CYGHWR_HAL_CORTEXM_STM32 == "F107VB") ||
                          (CYGHWR_HAL_CORTEXM_STM32 == "F107RC") || (CYGHWR_HAL_CORTEXM_STM32 == "F107VC") ||
			  (CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F2") ||
			  (CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F4") ||
			  (CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F7" )
                        }
        description     "Indicates that this part belongs to the connectivity
                         family of devices. These have slightly different interrupt
                         and GPIO layouts to the original STM32 F103 devices."
    }

    cdl_option CYGNUM_HAL_CORTEXM_PRIORITY_LEVEL_BITS {
        display         "CPU priority levels"
        flavor          data
        calculated      4
        description     "This option defines the number of bits used to
                         encode the exception priority levels that this
                         variant of the Cortex-M CPU implements."
    }

    cdl_component CYGHWR_HAL_CORTEXM_STM32_CLOCK {
        display         "Clock setup calculations"
        flavor          none
        no_define
        cdl_option CYGHWR_HAL_CORTEXM_STM32_CLOCK_PLL_SOURCE {
            display         "PLL input source"
            flavor          data
            default_value   { "HSE" }
            legal_values    { "HSI" "HSE" }
            description     "
                This sets whether the PLL will be driven by the external
                high-speed clock (HSE), or internal high-speed clock (HSI)."
        }

        cdl_option CYGHWR_HAL_CORTEXM_STM32_CLOCK_PLL_PREDIV {
            display         "PLL pre-divider"
            flavor          data
            default_value   1
            legal_values    1 to 63
            requires        { !CYGHWR_HAL_CORTEXM_STM32_CONNECTIVITY implies (CYGHWR_HAL_CORTEXM_STM32_CLOCK_PLL_PREDIV <= 2) }
            requires        { (CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F1") implies (CYGHWR_HAL_CORTEXM_STM32_CLOCK_PLL_PREDIV <= 16) }
            requires        { ((CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F1") && (CYGHWR_HAL_CORTEXM_STM32_CLOCK_PLL_SOURCE == "HSI")) implies \
                                  (CYGHWR_HAL_CORTEXM_STM32_CLOCK_PLL_PREDIV == 2) }
            requires        { ((CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F2") || (CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F4")) implies (CYGHWR_HAL_CORTEXM_STM32_CLOCK_PLL_PREDIV >= 2) }
	    requires        { (CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F7") implies (CYGHWR_HAL_CORTEXM_STM32_CLOCK_PLL_PREDIV >= 2) }
            description     "
               This option corresponds to the divider used before input to the PLL.
               On non-connectivity parts, you can only divide by 2 or 1. On other
               F1 parts, if using HSI as the clock source, then that is automatically
               divided by 2. If using HSE as the clock source, then this value corresponds
               to the PREDIV1 field of register RCC_CFGR2. On F2 and F4 parts, this value
               corresponds to the PLLM field of RCC_PLLCFGR."
        }


        cdl_option CYGHWR_HAL_CORTEXM_STM32_CLOCK_PLL_MUL {
            display         "PLL multiplier"
            flavor          data
            default_value   9
            legal_values    2 to 432
            requires        { (CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F1") implies (CYGHWR_HAL_CORTEXM_STM32_CLOCK_PLL_MUL <= 16) }
            requires        { ((CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F2") || (CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F4")) implies (CYGHWR_HAL_CORTEXM_STM32_CLOCK_PLL_MUL <= 432) }
            requires        { (CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F7") implies (CYGHWR_HAL_CORTEXM_STM32_CLOCK_PLL_MUL <= 432) }
            description     "
                This value is used to multiply up the PLL input. On the F1 it corresponds
                to the PLLMUL field of RCC_CFGR. On the F2 and F4 it corresponds to the PLLN
                field of RCC_PLLCFGR."
        }

        cdl_option CYGHWR_HAL_CORTEXM_STM32_CLOCK_SYSCLK_DIV {
            display         "SYSCLK divider"
            flavor          data
	    active_if       { ((CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F2") || (CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F4") || (CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F7")) }
            default_value   2
            legal_values    { 2 4 6 8 }
            description     "
                This value is used to divide down the PLL output for use as
                the SYSCLK clock. This corresponds to the PLLP field of
                RCC_PLLCFGR"
        }

        cdl_option CYGHWR_HAL_CORTEXM_STM32_CLOCK_HCLK_DIV {
            display         "HCLK divider"
            flavor          data
            default_value   1
            legal_values    { 1 2 4 8 16 64 128 256 512 }
            description     "Divider for AHB"
        }

        cdl_option CYGHWR_HAL_CORTEXM_STM32_CLOCK_PCLK1_DIV {
            display         "PCLK1 divider"
            flavor          data
            default_value   2
            legal_values    { 1 2 4 8 16 }
            description     "Divider for APB1"
        }

        cdl_option CYGHWR_HAL_CORTEXM_STM32_CLOCK_PCLK2_DIV {
            display         "PCLK2 divider"
            flavor          data
            default_value   1
            legal_values    { 1 2 4 8 16 }
            description     "Divider for APB2"
        }

        cdl_option CYGHWR_HAL_CORTEXM_STM32_CLOCK_PLLQ_DIV {
            display         "PLLQ divider"
            flavor          data
	    active_if       { ((CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F2") || (CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F4") || (CYGHWR_HAL_CORTEXM_STM32_FAMILY=="F7")) }
            default_value   7
            legal_values    4 to 15
            description     "
               This PLL divider is used in the F2 and F4 families to divide down the
               PLL output clock (VCO clock) for use by the USB OTG FS, SDIO
               and RNG peripherals. USB OTG FS requires a 48MHz clock and
               other peripherals require a clock no greater than 48MHz."
        }
    }

    cdl_option CYGNUM_HAL_KERNEL_COUNTERS_CLOCK_ISR_DEFAULT_PRIORITY {
        display       "Clock interrupt ISR priority"
        flavor        data
        calculated    0xE0
        description   "Set clock ISR priority to lowest priority."
    }

    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
        no_define
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            default_value 1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            default_value 1000000 / CYGNUM_HAL_RTC_DENOMINATOR
            description   "The period defined here is something of a fake, it is expressed
                           in terms of a notional 1MHz clock. The value actually installed
                           in the hardware is calculated from the current settings of the
                           clock generation hardware."
        }
    }

    cdl_interface CYGINT_HAL_STM32_UART0 {
        display     "Platform has UART0 serial port"
        description "The platform has a socket on UART0."
    }

    cdl_interface CYGINT_HAL_STM32_UART1 {
        display     "Platform has UART1 serial port"
        description "The platform has a socket on UART1."
    }

    cdl_interface CYGINT_HAL_STM32_UART2 {
        display     "Platform has UART2 serial port"
        description "The platform has a socket on UART2."
    }

    cdl_interface CYGINT_HAL_STM32_UART3 {
        display     "Platform has UART3 serial port"
        description "The platform has a socket on UART3."
    }

    cdl_interface CYGINT_HAL_STM32_UART4 {
        display     "Platform has UART4 serial port"
        description "The platform has a socket on UART4."
    }

    cdl_interface CYGINT_HAL_STM32_UART5 {
        display     "Platform has UART5 serial port"
        description "The platform has a socket on UART5."
    }

    cdl_component CYGHWR_HAL_STM32_UART0_REMAP {
        display       "Remap UART0 (USART1) pins"
	flavor	      bool
        default_value 0

        description   "Remap UART0 (USART1) to alternate set of pins.
                       This will usually be set by the platform
                       HAL to reflect the configuration of the hardware."

	cdl_option CYGHWR_HAL_STM32_UART0_PIN_TX {
	    display       "TX pin"
	    active_if	  (CYGHWR_HAL_STM32_UART0_REMAP == 1)
	    flavor        data
	    default_value { "A, 9" }
	    legal_values  { "A, 9" "B, 6" }

	    description   "This option specifies the pin of TX serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART0_PIN_RX {
	    display       "RX pin"
	    active_if	  (CYGHWR_HAL_STM32_UART0_REMAP == 1)
	    flavor        data
	    default_value { "A, 10" }
	    legal_values  { "A, 10" "B, 7" }

	    description   "This option specifies the pin of RX serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART0_PIN_CTS {
	    display       "CTS pin"
	    active_if	  (CYGHWR_HAL_STM32_UART0_REMAP == 1)
	    flavor        data
	    default_value { "A, 11" }
	    legal_values  { "A, 11" }

	    description   "This option specifies the pin of CTS serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART0_PIN_RTS {
	    display       "RTS pin"
	    active_if	  (CYGHWR_HAL_STM32_UART0_REMAP == 1)
	    flavor        data
	    default_value { "A, 12" }
	    legal_values  { "A, 12" }

	    description   "This option specifies the pin of RTS serial device."
	}
    }

    cdl_component CYGHWR_HAL_STM32_UART1_REMAP {
        display       "Remap UART1 (USART2) pins"
	flavor	      bool
        default_value 0

        description   "Remap UART1 (USART2) to alternate set of pins.
                       This will usually be set by the platform
                       HAL to reflect the configuration of the hardware."

	cdl_option CYGHWR_HAL_STM32_UART1_PIN_TX {
	    display       "TX pin"
	    active_if	  (CYGHWR_HAL_STM32_UART1_REMAP == 1)
	    flavor        data
	    default_value { "A, 2" }
	    legal_values  { "A, 2" "D, 5" }

	    description   "This option specifies the pin of TX serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART1_PIN_RX {
	    display       "RX pin"
	    active_if	  (CYGHWR_HAL_STM32_UART1_REMAP == 1)
	    flavor        data
	    default_value { "A, 3" }
	    legal_values  { "A, 3" "D, 6" }

	    description   "This option specifies the pin of RX serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART1_PIN_CTS {
	    display       "CTS pin"
	    active_if	  (CYGHWR_HAL_STM32_UART1_REMAP == 1)
	    flavor        data
	    default_value { "A, 0" }
	    legal_values  { "A, 0" "D, 3" }

	    description   "This option specifies the pin of CTS serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART1_PIN_RTS {
	    display       "RTS pin"
	    active_if	  (CYGHWR_HAL_STM32_UART1_REMAP == 1)
	    flavor        data
	    default_value { "A, 1" }
	    legal_values  { "A, 1" "D, 4" }

	    description   "This option specifies the pin of RTS serial device."
	}
    }

    # CYGHWR_HAL_CORTEXM_STM32_FAMILY_F1 left for
    # backward compatibility with familiy F1
    # New remap was added with _N suffix in contradiction to
    # other REMAPs
    cdl_option CYGHWR_HAL_STM32_UART2_REMAP {
        display       "Remap UART2 (USART3) pins"
	active_if     { CYGHWR_HAL_CORTEXM_STM32_FAMILY_F1 }
	flavor	      data
        default_value { "NONE" }
        legal_values  { "NONE" "PARTIAL" "FULL" }

        description   "Remap UART2 (USART3) to alternate set of pins.
                       This will usually be set by the platform
                       HAL to reflect the configuration of the hardware."
    }

    cdl_component CYGHWR_HAL_STM32_UART2_REMAP_N {
        display       "Remap UART2 (USART3) pins"
	active_if     { !CYGHWR_HAL_CORTEXM_STM32_FAMILY_F1 }
	flavor	      bool
        default_value 0

        description   "Remap UART2 (USART3) to alternate set of pins.
                       This will usually be set by the platform
                       HAL to reflect the configuration of the hardware."

	cdl_option CYGHWR_HAL_STM32_UART2_PIN_TX {
	    display       "TX pin"
	    active_if	  (CYGHWR_HAL_STM32_UART2_REMAP_N == 1)
	    flavor        data
	    default_value { "B, 10" }
	    legal_values  { "B, 10" "D, 8" "C, 10" }

	    description   "This option specifies the pin of TX serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART2_PIN_RX {
	    display       "RX pin"
	    active_if	  (CYGHWR_HAL_STM32_UART2_REMAP_N == 1)
	    flavor        data
	    default_value { "B, 11" }
	    legal_values  { "B, 11" "D, 9" "C, 11" }

	    description   "This option specifies the pin of RX serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART2_PIN_CTS {
	    display       "CTS pin"
	    active_if	  (CYGHWR_HAL_STM32_UART2_REMAP_N == 1)
	    flavor        data
	    default_value { "B, 13" }
	    legal_values  { "B, 13" "D, 11" }

	    description   "This option specifies the pin of CTS serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART2_PIN_RTS {
	    display       "RTS pin"
	    active_if	  (CYGHWR_HAL_STM32_UART2_REMAP_N == 1)
	    flavor        data
	    default_value { "B, 14" }
	    legal_values  { "B, 14" "D, 12" }

	    description   "This option specifies the pin of RTS serial device."
	}
    }

    cdl_component CYGHWR_HAL_STM32_UART3_REMAP {
        display       "Remap UART3 (UART4) pins"
	flavor	      bool
        default_value 0

        description   "Remap UART3 (UART4) to alternate set of pins.
                       This will usually be set by the platform
                       HAL to reflect the configuration of the hardware."

	cdl_option CYGHWR_HAL_STM32_UART3_PIN_TX {
	    display       "TX pin"
	    active_if	  (CYGHWR_HAL_STM32_UART3_REMAP == 1)
	    flavor        data
	    requires	  { CYGHWR_HAL_STM32_UART1_PIN_CTS != CYGHWR_HAL_STM32_UART3_PIN_TX }
	    requires	  { CYGHWR_HAL_STM32_UART2_PIN_TX  != CYGHWR_HAL_STM32_UART3_PIN_TX }
	    default_value { "A, 0" }
	    legal_values  { "A, 0" "C, 10" }

	    description   "This option specifies the pin of TX serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART3_PIN_RX {
	    display       "RX pin"
	    active_if	  (CYGHWR_HAL_STM32_UART3_REMAP == 1)
	    flavor        data
	    requires	  { CYGHWR_HAL_STM32_UART1_PIN_RTS != CYGHWR_HAL_STM32_UART3_PIN_RX }
	    requires	  { CYGHWR_HAL_STM32_UART2_PIN_RX  != CYGHWR_HAL_STM32_UART3_PIN_RX }
	    default_value { "A, 1" }
	    legal_values  { "A, 1" "C, 11" }

	    description   "This option specifies the pin of RX serial device."
	}
    }

    cdl_component CYGHWR_HAL_STM32_UART4_REMAP {
        display       "Remap UART4 (UART5) pins"
	flavor	      bool
        default_value 0

        description   "Remap UART4 (UART5) to alternate set of pins.
                       This will usually be set by the platform
                       HAL to reflect the configuration of the hardware."

	cdl_option CYGHWR_HAL_STM32_UART4_PIN_TX {
	    display       "TX pin"
	    active_if	  (CYGHWR_HAL_STM32_UART4_REMAP == 1)
	    flavor        data
	    default_value { "C, 12" }
	    legal_values  { "C, 12" }

	    description   "This option specifies the pin of TX serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART4_PIN_RX {
	    display       "RX pin"
	    active_if	  (CYGHWR_HAL_STM32_UART4_REMAP == 1)
	    flavor        data
	    default_value { "D, 2" }
	    legal_values  { "D, 2" }

	    description   "This option specifies the pin of RX serial device."
	}
    }

    cdl_component CYGHWR_HAL_STM32_UART5_REMAP {
        display       "Remap UART5 (USART6) pins"
	flavor	      bool
        default_value 0

        description   "Remap UART5 (USART6) to alternate set of pins.
                       This will usually be set by the platform
                       HAL to reflect the configuration of the hardware."

	cdl_option CYGHWR_HAL_STM32_UART5_PIN_TX {
	    display       "TX pin"
	    active_if	  (CYGHWR_HAL_STM32_UART5_REMAP == 1)
	    flavor        data
	    default_value { "C, 6" }
	    legal_values  { "C, 6" "G, 14" }

	    description   "This option specifies the pin of TX serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART5_PIN_RX {
	    display       "RX pin"
	    active_if	  (CYGHWR_HAL_STM32_UART5_REMAP == 1)
	    flavor        data
	    default_value { "C, 7" }
	    legal_values  { "C, 7" "G, 9" }

	    description   "This option specifies the pin of RX serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART5_PIN_CTS {
	    display       "CTS pin"
	    active_if	  (CYGHWR_HAL_STM32_UART5_REMAP == 1)
	    flavor        data
	    default_value { "G, 13" }
	    legal_values  { "G, 13" "G, 15" }

	    description   "This option specifies the pin of CTS serial device."
	}

	cdl_option CYGHWR_HAL_STM32_UART5_PIN_RTS {
	    display       "RTS pin"
	    active_if	  (CYGHWR_HAL_STM32_UART5_REMAP == 1)
	    flavor        data
	    default_value { "G, 8" }
	    legal_values  { "G, 8" "G, 12" }

	    description   "This option specifies the pin of RTS serial device."
	}
    }

    cdl_component CYGHWR_HAL_STM32_I2C1_REMAP {
        display       "Remap I2C bus 1 pins"
        flavor        bool
        default_value 0

        description   "Remap I2C bus 1 to alternate set of pins."

	    cdl_option CYGHWR_HAL_STM32_I2C1_SDA {
		display		"SDA"
		active_if	(CYGHWR_HAL_STM32_I2C1_REMAP == 1)
		flavor		data
		default_value	{ "B, 9" }
		legal_values	{ "B, 9" "B, 7" }
		description "
		    This option specifies the SDA pin."
	    }

	    cdl_option CYGHWR_HAL_STM32_I2C1_SCL {
		display		"SCL"
		active_if	(CYGHWR_HAL_STM32_I2C1_REMAP == 1)
		flavor		data
		default_value	{ "B, 8" }
		legal_values	{ "B, 8" "B, 6" }
		description "
		    This option specifies the SCL pin."
	    }
    }

    cdl_component CYGHWR_HAL_STM32_I2C2_REMAP {
        display       "Remap I2C bus 2 pins"
        flavor        bool
        default_value 0

        description   "Remap I2C bus 2 to alternate set of pins."

	    cdl_option CYGHWR_HAL_STM32_I2C2_SDA {
		display		"SDA"
		active_if	(CYGHWR_HAL_STM32_I2C2_REMAP == 1)
		flavor		data
		default_value	{ "B, 11" }
		legal_values	{ "B, 11" "F, 0" "H, 5" }
		description	"This option specifies the SDA pin."
	    }

	    cdl_option CYGHWR_HAL_STM32_I2C2_SCL {
		display		"SCL"
		active_if	(CYGHWR_HAL_STM32_I2C2_REMAP == 1)
		flavor		data
		default_value	{ "B, 10" }
		legal_values	{ "B, 10" "F, 1" "H, 4" }
		description	"This option specifies the SCL pin."
	    }
    }

    cdl_component CYGHWR_HAL_STM32_I2C3_REMAP {
        display       "Remap I2C bus 3 pins"
	flavor	      bool
        default_value 0

        description   "Remap I2C bus 3 to alternate set of pins."

	    cdl_option CYGHWR_HAL_STM32_I2C3_SDA {
		display		"SDA"
		active_if	(CYGHWR_HAL_STM32_I2C3_REMAP == 1)
		flavor		data
		default_value	{ "C, 9" }
		legal_values	{ "C, 9" "H, 8" }
		description	"This option specifies the SDA pin."
	    }

	    cdl_option CYGHWR_HAL_STM32_I2C3_SCL {
		display		"SCL"
		active_if	(CYGHWR_HAL_STM32_I2C3_REMAP == 1)
		flavor		data
		default_value	{ "A, 8" }
		legal_values	{ "A, 8" "H, 7" }
		description	"This option specifies the SCL pin."
	    }
    }

    cdl_component CYGHWR_HAL_STM32_SPI1_REMAP {
        display       "Remap SPI bus 1 pins"
        active_if     CYGHWR_HAL_CORTEXM_STM32_CONNECTIVITY
        flavor        bool
        default_value 0

        description   "Remap SPI bus 1 to alternate set of pins.
		       This option is only available on connectivity line
                       devices."

		cdl_option CYGHWR_HAL_STM32_SPI1_PIN_MOSI {
			display       "MOSI pin"
			active_if     (CYGHWR_HAL_STM32_SPI1_REMAP == 1)
			flavor        data
			default_value { "A, 7" }
			legal_values  { "A, 7" "B, 5" }

			description   "This option specifies the pin of MOSI."
		}

		cdl_option CYGHWR_HAL_STM32_SPI1_PIN_MISO {
			display       "MISO pin"
			active_if     (CYGHWR_HAL_STM32_SPI1_REMAP == 1)
			flavor        data
			default_value { "A, 6" }
			legal_values  { "A, 6" "B, 4" }

			description   "This option specifies the pin of MISO."
		}

		cdl_option CYGHWR_HAL_STM32_SPI1_PIN_SCK {
			display       "SCK pin"
			active_if     (CYGHWR_HAL_STM32_SPI1_REMAP == 1)
			flavor        data
			default_value { "A, 5" }
			legal_values  { "A, 5" "B, 3" }

			description   "This option specifies the pin of SCK."
		}

		cdl_option CYGHWR_HAL_STM32_SPI1_PUPD {
			display       "PUPD out resistor"
			active_if     (CYGHWR_HAL_STM32_SPI1_REMAP == 1)
			flavor        data
			default_value { "NONE" }
			legal_values  { "NONE" "PULLUP" "PULLDOWN" }

			description   "This option specifies the PUPD mode."
		}
    }

    cdl_component CYGHWR_HAL_STM32_SPI2_REMAP {
        display       "Remap SPI bus 2 pins"
        active_if     CYGHWR_HAL_CORTEXM_STM32_CONNECTIVITY
        flavor        bool
        default_value 0

        description   "Remap SPI bus 2 to alternate set of pins.
		       This option is only available on connectivity line
                       devices."

		cdl_option CYGHWR_HAL_STM32_SPI2_PIN_MOSI {
			display       "MOSI pin"
			active_if     (CYGHWR_HAL_STM32_SPI2_REMAP == 1)
			flavor        data
			default_value { "B, 15" }
			legal_values  { "B, 15" "C, 3" "I, 3" }

			description   "This option specifies the pin of MOSI."
		}

		cdl_option CYGHWR_HAL_STM32_SPI2_PIN_MISO {
			display       "MISO pin"
			active_if     (CYGHWR_HAL_STM32_SPI2_REMAP == 1)
			flavor        data
			default_value { "B, 14" }
			legal_values  { "B, 14" "C, 2" "I, 2" }

			description   "This option specifies the pin of MISO."
		}

		cdl_option CYGHWR_HAL_STM32_SPI2_PIN_SCK {
			display       "SCK pin"
			active_if     (CYGHWR_HAL_STM32_SPI2_REMAP == 1)
			flavor        data
			default_value { "B, 13" }
			legal_values  { "B, 10" "B, 13" "D, 3" "I, 1" }

			description   "This option specifies the pin of SCK."
		}

		cdl_option CYGHWR_HAL_STM32_SPI2_PUPD {
			display       "PUPD out resistor"
			active_if     (CYGHWR_HAL_STM32_SPI2_REMAP == 1)
			flavor        data
			default_value { "NONE" }
			legal_values  { "NONE" "PULLUP" "PULLDOWN" }

			description   "This option specifies the PUPD mode."
		}
    }

    cdl_component CYGHWR_HAL_STM32_SPI3_REMAP {
        display       "Remap SPI bus 3 pins"
        active_if     CYGHWR_HAL_CORTEXM_STM32_CONNECTIVITY
        flavor        bool
        default_value 0

        description   "Remap SPI bus 3 to alternate set of pins.
                       This option is only available on connectivity line
                       devices."

		cdl_option CYGHWR_HAL_STM32_SPI3_PIN_MOSI {
			display       "MOSI pin"
			active_if     (CYGHWR_HAL_STM32_SPI3_REMAP == 1)
			flavor        data
			default_value { "B, 5" }
			legal_values  { "B, 5" "C, 12" "D, 6" }

			description   "This option specifies the pin of MOSI."
		}

		cdl_option CYGHWR_HAL_STM32_SPI3_PIN_MISO {
			display       "MISO pin"
			active_if     (CYGHWR_HAL_STM32_SPI3_REMAP == 1)
			flavor        data
			default_value { "B, 4" }
			legal_values  { "B, 4" "C, 11" }

			description   "This option specifies the pin of MISO."
		}

		cdl_option CYGHWR_HAL_STM32_SPI3_PIN_SCK {
			display       "SCK pin"
			active_if     (CYGHWR_HAL_STM32_SPI3_REMAP == 1)
			flavor        data
			default_value { "B, 3" }
			legal_values  { "B, 3" "C, 10" }

			description   "This option specifies the pin of SCK."
		}

		cdl_option CYGHWR_HAL_STM32_SPI3_PUPD {
			display       "PUPD out resistor"
			active_if     (CYGHWR_HAL_STM32_SPI3_REMAP == 1)
			flavor        data
			default_value { "NONE" }
			legal_values  { "NONE" "PULLUP" "PULLDOWN" }

			description   "This option specifies the PUPD mode."
		}

		cdl_option CYGHWR_HAL_STM32_SPI3_MOSI_DAF {
			display       "MOSI AF register"
			active_if     ( CYGHWR_HAL_STM32_SPI3_REMAP == 1)
			calculated    { CYGHWR_HAL_STM32_SPI3_PIN_MOSI == "D, 6" ? 1 : 0 }

			description   "This option specifies AF register for MOSI."
		}
    }

    cdl_component CYGHWR_HAL_STM32_SPI5_REMAP {
        display       "Remap SPI bus 5 pins"
        active_if     CYGHWR_HAL_CORTEXM_STM32_CONNECTIVITY
        flavor        bool
        default_value 0

        description   "Remap SPI bus 5 to alternate set of pins.
                       This option is only available on connectivity line
                       devices."

		cdl_option CYGHWR_HAL_STM32_SPI5_PIN_MOSI {
			display       "MOSI pin"
			active_if     (CYGHWR_HAL_STM32_SPI5_REMAP == 1)
			flavor        data
			default_value { "F, 9" }
			legal_values  { "F, 9" "F, 11" }

			description   "This option specifies the pin of MOSI."
		}

		cdl_option CYGHWR_HAL_STM32_SPI5_PIN_MISO {
			display       "MISO pin"
			active_if     (CYGHWR_HAL_STM32_SPI5_REMAP == 1)
			flavor        data
			default_value { "F, 8" }
			legal_values  { "F, 8" "H, 7" }

			description   "This option specifies the pin of MISO."
		}

		cdl_option CYGHWR_HAL_STM32_SPI5_PIN_SCK {
			display       "SCK pin"
			active_if     (CYGHWR_HAL_STM32_SPI5_REMAP == 1)
			flavor        data
			default_value { "F, 7" }
			legal_values  { "F, 7" "H, 6" }

			description   "This option specifies the pin of SCK."
		}

		cdl_option CYGHWR_HAL_STM32_SPI5_PUPD {
			display       "PUPD out resistor"
			active_if     (CYGHWR_HAL_STM32_SPI5_REMAP == 1)
			flavor        data
			default_value { "NONE" }
			legal_values  { "NONE" "PULLUP" "PULLDOWN" }

			description   "This option specifies the PUPD mode."
		}
    }

    cdl_option CYGFUN_HAL_CORTEXM_STM32_PROFILE_TIMER {
        display       "Use TIM2 for gprof profiling"
        active_if     CYGPKG_PROFILE_GPROF
        flavor        bool
        default_value 1
        implements    CYGINT_PROFILE_HAL_TIMER
        implements    CYGINT_HAL_COMMON_SAVED_INTERRUPT_STATE_REQUIRED
        description   "
            The STM32 variant HAL can provide support for gprof-based
            profiling. This uses timer TIM2 to generate regular interrupts,
            and the interrupt handler records the PC at the time of the
            interrupt. Disable this option if you wish to provide
            an alternative profiling timer implementation."
    }

    cdl_component CYGPKG_HAL_CORTEXM_STM32_OPTIONS {
        display "Build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package."

        cdl_option CYGPKG_HAL_CORTEXM_STM32_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the STM32 variant HAL package. These flags are used
                in addition to the set of global flags."
        }

        cdl_option CYGPKG_HAL_CORTEXM_STM32_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the STM32 variant HAL package. These flags are removed from
                the set of global flags if present."
        }
    }

    cdl_option CYGPKG_HAL_CORTEXM_STM32_TESTS {
        display "STM32 tests"
        active_if      CYGPKG_KERNEL
        flavor  data
        no_define
        calculated { "tests/timers" }
        description   "
            This option specifies the set of tests for the STM32 HAL."
    }
}

# EOF hal_cortexm_stm32.cdl
