# ====================================================================
#
#      olpce2294_eth_drivers.cdl
#
#      Ethernet drivers - platform dependent support for OLPCE2294
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2008 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Sergei Gavrikov
# Contributors:   Sergei Gavrikov
# Date:           2008-08-31
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_ARM_OLPCE2294 {
    display       "LAN ethernet driver for Olimex LPC-E2294"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_HAL_ARM_LPC2XXX_OLPCE2294

    implements    CYGINT_DEVS_ETH_CL_CS8900A_REQUIRED

    requires      CYGPKG_DEVS_ETH_CL_CS8900A

    # Olimex LPC-E2294 development board has Cirrus Logic CS8900A ethernet
    # controller had been wired in a dumb 8-bit mode.
    requires      CYGIMP_DEVS_ETH_CL_CS8900A_DATABUS_8BIT

    include_dir   cyg/io

    description   "
        Ethernet driver for Olimex LPC-E2294 board."

    cdl_interface CYGINT_DEVS_ETH_CL_CS8900A_REQUIRED {
        display   "CL CS8900A ethernet driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_CL_CS8900A_INL <cyg/io/devs_eth_arm_olpce2294.inl>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_CL_CS8900A_CFG <pkgconf/devs_eth_arm_olpce2294.h>"
        puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
    }

    cdl_component CYGSEM_DEVS_ETH_CL_CS8900A_NOINTS {
        display       "Interrupts are not supported"
        calculated    1
        description   "
            Interrups are not supported in 8-bit mode. Polled mode must
            be used."
    }

   cdl_component CYGPKG_DEVS_ETH_ARM_OLPCE2294_ETH0 {
        display       "OLPCE2294 ethernet port driver"
        flavor        bool
        default_value 1
        description   "
            This option includes the ethernet device driver for the
            OLPCE2294 port."

        implements CYGHWR_NET_DRIVER_ETH0
        implements CYGINT_DEVS_ETH_CL_CS8900A_REQUIRED
        implements CYGINT_DEVS_ETH_CL_CS8900A_DATABUS_8BIT

        cdl_option CYGDAT_DEVS_ETH_ARM_OLPCE2294_ETH0_NAME {
            display       "Device name for the ETH0 ethernet driver"
            flavor        data
            default_value {"\"eth0\""}
            description   "
                This option sets the name of the ethernet device."
        }

	cdl_component CYGSEM_DEVS_ETH_ARM_OLPCE2294_ETH0_SET_ESA {
	    display       "Set the ethernet station address"
	    flavor        bool
	    calculated    1
	    description   "Enabling this option will allow the ethernet
	    station address to be forced to the value set by the
	    configuration."

	    cdl_option CYGDAT_DEVS_ETH_ARM_OLPCE2294_ETH0_ESA {
	        display       "The ethernet station address"
	        flavor        data
	        default_value {"{0x08, 0x88, 0x12, 0x34, 0x56, 0x78}"}
	        description   "The ethernet station address"
	    }
	}
    }
}

