# ====================================================================
#
#      cl_cs8900a_eth_drivers.cdl
#
#      Ethernet driver for Cirrus Logic CS8900A controller
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Contributors:   gthomas, jskov
# Date:           2001-11-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_CL_CS8900A {
    display       "Driver for Cirrus Logic CS8900A ethernet controller."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS

    implements    CYGHWR_NET_DRIVERS
    implements    CYGINT_IO_ETH_MULTICAST

    active_if     CYGINT_DEVS_ETH_CL_CS8900A_REQUIRED

    include_dir   cyg/io
    description   "Driver for Cirrus Logic CS8900A ethernet controller."
    compile       -library=libextras.a if_cs8900a.c

    define_proc {
        puts $::cdl_header "#include <pkgconf/system.h>";
        puts $::cdl_header "#include CYGDAT_DEVS_ETH_CL_CS8900A_CFG";
    }

    cdl_option CYGSEM_DEVS_ETH_CL_CS8900A_WRITE_EEPROM {
        display "SIOCSIFHWADDR records ESA (MAC address) in EEPROM"
        default_value 0
        description   "
            The ioctl() socket call with operand SIOCSIFHWADDR sets the
            interface hardware address - the MAC address or Ethernet Station
            Address (ESA).  This option causes the new MAC address to be written
            into the EEPROM associated with the interface, so that the new
            MAC address is permanently recorded.  Doing this should be a
            carefully chosen decision, hence this option."
    }

    cdl_option CYGIMP_DEVS_ETH_CL_CS8900A_DATABUS_8BIT {
        display "8-bit data bus"
        flavor        bool
        requires      !CYGSEM_DEVS_ETH_CL_CS8900A_WRITE_EEPROM
        requires      CYGSEM_DEVS_ETH_CL_CS8900A_NOINTS
        default_value 0
        description   "
            The CS8900A can been use in 8-bit mode. From AN181 from
            Cirrus Logic... Unsupported functions in 8-bit mode:
            Interrupts are not supported. Polled mode must be used;
            The DMA engine only uses 16 bit memory access and does not
            support 8 bit transfers; The packet page pointer has an
            auto increment feature that cannot be used in 8-bit mode;
            An EEPROM is not supported."
    }

    cdl_option CYGIMP_DEVS_ETH_CL_CS8900A_DATABUS_BYTE_SWAPPED {
	display "Byte swapped data bus"
	flavor  bool
	default_value 0
	description   "
		    From the application note AN205 from Cirrus Logic ...The CS8900a
			assumes a litte-endian ISA type system. However, network byte order
			is always big-endian.Therefore to minimize software manipulation of
			frame data in ISA systems, the CS8900 byte-swaps frame data
			internally. The control and status registers are not byte-swapped.
			In a big-endian system you can either byte-swap the network data
			(to reverse the byte swapping done internally to the CS8900) in
			software or you can do it in hardware (byte swap the data lines to
			the chip). Byte swapping the data lines is much more efficient; you
	        will only need to byte swap the control/status/counter values in
			software and not the frame data. (Most of the read/writes to the chip
			are frame data.) Since network byte order is always big endian, this
		    scheme works without special support on the other end of the network...
			Normally, you won't need to check this option unless you are using a
			CS8900a ethernet controller with a big endian machine and hardware
			that has been designed with the cs8900a in mind."
    }

    cdl_component CYGPKG_DEVS_ETH_CL_CS8900A_OPTIONS {
        display "Cirrus Logic ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_CL_CS8900A_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the Cirrus Logic ethernet driver package.
                These flags are used in addition
                to the set of global flags."
        }
    }
}

