# ====================================================================
#
#      i2c_lpc2xxx.cdl
#
#      eCos LPC2xxx I2C configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Hans Rosenfeld <rosenfeld@grumpf.hope-2000.org>
# Contributors:   Uwe Kindler <uwe_kindler@web.de>
# Date:           2007-07-12
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_I2C_ARM_LPC2XXX {
    display     "I2C driver for LPC2xxx family of ARM controllers"
    
    parent      CYGPKG_IO_I2C
    active_if   CYGPKG_IO_I2C
    active_if   CYGPKG_HAL_ARM_LPC2XXX || CYGPKG_HAL_ARM_LPC24XX 

    description " 
           This package provides a generic I2C device driver for the on-chip
           I2C peripherals in LPX2xxx processors."
           
    include_dir cyg/io
    compile     i2c_lpc2xxx.c
    
    cdl_option CYGHWR_DEVS_I2C_ARM_LPC2XXX_MULTIPLE_BUSES {
	display		"Target hardware may have multiple I2C buses"
	flavor		bool
	default_value	0
	description "
          The LPC2xxx I2C driver can support multiple I2C bus devices. By
          default the driver assumes only a single device is present and will
          optimize for that case, using constant definitions provided by the
          platform HAL rather than per-device structure fields. If the hardware
          has multiple I2C bus devices, or if a singleton bus is instantiated
          by some other package and hence the platform HAL cannot provide the
          necessary definitions, then this option should be enabled."
    }
    
    cdl_option CYGPKG_DEVS_I2C_ARM_LPC2XXX_DEBUG_LEVEL {
         display "Driver debug output level"
         flavor  data
         legal_values {0 1}
         default_value 0
         description   "
             This option specifies the level of debug data output by
             the LPC2XXX I2C device driver. A value of 0 signifies
             no debug data output; 1 signifies normal debug data
             output. The generic eCos I2C driver functions do not return any 
             error information if a I2C transfer failed. If this option is
             1 then the driver prints the status flags if a transfer failed
             or was aborted. It prints the status flags in case of a missing 
             data or address acknowledge, in case of lost arbitration and in 
             case of a bus error. A missing acknowledge does not realy indicate
             an error and may be part of a normal I2C communication. Therefore
             this option should only be >0 for debug reasons."         
    }
}
