##==========================================================================
##
##      hal_freescale_edma.cdl
##
##      Cortex-M Freescale Kinetis eDMA
##
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##==========================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):    Ilija Kocho <ilijak@siva.com.mk>
## Date:         2011-12-11
##
######DESCRIPTIONEND####
##
##==========================================================================

cdl_package CYGPKG_HAL_FREESCALE_EDMA {
    display "Freescale eDMA controller"
    hardware

    include_dir cyg/hal
    compile hal_freescale_edma.c
    
    active_if CYGINT_HAL_DMA

    cdl_option CYGNUM_HAL_FREESCALE_EDMA_CHAN_NUM {
        display "Number of DMA channels"
        flavor data
        legal_values { 16 32 }
        default_value 16
    }

    cdl_option CYGOPT_HAL_FREESCALE_EDMA_ERCA {
        display "Round robin channel arbitration"
        flavor bool
        default_value 0
    }

    cdl_option CYGOPT_HAL_FREESCALE_EDMA_EMLM {
        display "Enable minor loop mapping"
        flavor bool
        default_value 1
    }

    cdl_option CYGOPT_HAL_FREESCALE_EDMA_CLM {
        display "Continuous link mode"
        flavor bool
        active_if CYGOPT_HAL_FREESCALE_EDMA_EMLM
        default_value 0
    }

    cdl_option CYGNUM_HAL_FREESCALE_EDMA_GROUP_SIZE {
        display "Number of channels in DMA group"
        flavor data
        calculated  16
    }

    cdl_component CYGHWR_HAL_FREESCALE_EDMA_GROPS {
        display "Groups"
        flavor none
        no_define
        active_if { CYGNUM_HAL_FREESCALE_EDMA_CHAN_NUM >
            CYGNUM_HAL_FREESCALE_EDMA_GROUP_SIZE }

        cdl_option CYGNUM_HAL_FREESCALE_EDMA_GROUP_NUM {
            display "Number of DMA groups"
            flavor data
            calculated  { CYGNUM_HAL_FREESCALE_EDMA_GROUP_SIZE ?
                CYGNUM_HAL_FREESCALE_EDMA_CHAN_NUM /
                CYGNUM_HAL_FREESCALE_EDMA_GROUP_SIZE : 0}
        }

        cdl_option CYGNUM_HAL_FREESCALE_EDMA_GR0_PRIO {
            display "Group 0 priority"
            flavor data
            legal_values 0 1
            default_value 0
        }

        cdl_option CYGNUM_HAL_FREESCALE_EDMA_GR1_PRIO {
            display "Group 1 priority"
            flavor data
            legal_values 0 1
            calculated { CYGNUM_HAL_FREESCALE_EDMA_GR0_PRIO ? 0 : 1 }
        }

        cdl_option CYGOPT_HAL_FREESCALE_EDMA_ERGA {
            display "Round robin group arbitration"
            active_if { CYGNUM_HAL_FREESCALE_EDMA_GROUP_NUM > 1 }
            flavor bool
            default_value 0
        }
    }

    cdl_option CYGNUM_HAL_FREESCALE_DMAMUX_CHAN_NUM {
        display "Channels per DMAMUX"
        flavor data
        calculated 16
    }

    cdl_component CYGNUM_HAL_FREESCALE_DMAMUX_NUM {
        display "Number of DMAMUX units"
        flavor data
        active_if { CYGNUM_HAL_FREESCALE_EDMA_CHAN_NUM >
            CYGNUM_HAL_FREESCALE_DMAMUX_CHAN_NUM
        }
        calculated { CYGNUM_HAL_FREESCALE_DMAMUX_CHAN_NUM ?
           ( CYGNUM_HAL_FREESCALE_EDMA_CHAN_NUM /
            CYGNUM_HAL_FREESCALE_DMAMUX_CHAN_NUM ) : 0
        }
    }
}

# EOF hal_freescale_dma.cdl
