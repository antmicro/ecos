# ====================================================================
#
#      flash_sh_se77x9.cdl
#
#      FLASH memory - Hardware support on Hitachi SH/SE77X9
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  jskov
# Contributors:
# Date:           2001-05-28
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_SH_SE77X9 {
    display       "Hitachi SH/SE77X9 FLASH memory support"

    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH
    requires	  CYGPKG_HAL_SH_SH77X9_SE77X9

    compile       sh_se77x9_flash.c

    # Arguably this should do in the generic package
    # but then there is a logic loop so you can never enable it.
    cdl_interface CYGINT_DEVS_FLASH_AMD_AM29XXXXX_REQUIRED {
        display   "Generic AMD flash driver required"
    }

    implements    CYGINT_DEVS_FLASH_AMD_AM29XXXXX_REQUIRED
    requires      CYGHWR_DEVS_FLASH_AMD_AM29LV160
}
