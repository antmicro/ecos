# ====================================================================
#
#      hal_mips_sim.cdl
#
#      MIPS SIM HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  bartv
# Contributors:
# Date:           1999-11-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_MIPS_SIM {
    display  "Minimal simulator"
    parent        CYGPKG_HAL_MIPS
    define_header hal_mips_sim.h
    include_dir   cyg/hal
    description   "
           The minimal simulator HAL package is provided for when only
           a simple simulation of the processor architecture is
           desired, as opposed to detailed simulation of any specific
           board. To use this minimal simulator the command
           `target sim --board=jmr3904pal' should be used from inside
           gdb. It is not possible to use any of the eCos device
           drivers when the simulator is running in this mode"

    compile       hal_diag.c platform.S plf_misc.c

    implements CYGINT_HAL_DEBUG_GDB_CTRLC_UNSUPPORTED

    cdl_option CYGBLD_HAL_TARGET_H {
        display "architecture header file"
        flavor data
        no_define
	define -file system.h CYGBLD_HAL_TARGET_H
        calculated { CYGPKG_HAL_MIPS_TX39 ? "<pkgconf/hal_mips_tx39.h>" :
                                            "<pkgconf/hal_mips_vr4300.h>"}
    }

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_mips_sim.h>"
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM"}
        default_value {"RAM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
            Only supports RAM startup."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            default_value 1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
        }
        # Isn't a nice way to handle freq requirement!
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            default_value 999
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { CYGPKG_HAL_MIPS_TX39 ? "mips-tx39-elf" : \
						   "mips64vr4300-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGBLD_GLOBAL_WARNFLAGS .
                            (CYGPKG_HAL_MIPS_TX39 ? "" : "-mgp32 -EB") .
                            " -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions "
            }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { (CYGPKG_HAL_MIPS_TX39 ? "" : "-mgp32 -EB") . " -g -nostdlib -Wl,--gc-sections -Wl,-static" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYGPKG_HAL_MIPS_TX39 ? "mips_tx39_sim_ram" :
                                            "mips_vr4300_sim_ram" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYGPKG_HAL_MIPS_TX39 ? "<pkgconf/mlt_mips_tx39_sim_ram.ldi>" :
                                                "<pkgconf/mlt_mips_vr4300_sim_ram.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYGPKG_HAL_MIPS_TX39 ? "<pkgconf/mlt_mips_tx39_sim_ram.h>" : 
                                                "<pkgconf/mlt_mips_vr4300_sim_ram.h>" }
        }
    }
}
