##==========================================================================
##
##      hal_cortexm_kinetis_kwikstik.cdl
##
##      Cortex-M Freescale KwikStik platform HAL configuration data
##
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2011, 2012 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
##==========================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):    Tomas Frydrych <tomas@sleepfive.com>
## Contributor(s): jld
## Date:         2011-12-15
## Original:     hal_cortexm_kinetis_twr_k40x256.cdl by Ilija Kocho
##
######DESCRIPTIONEND####
##
##==========================================================================

cdl_package CYGPKG_HAL_CORTEXM_KINETIS_KWIKSTIK {
    display       "Freescale Kinetis KwikStik Platform"
    parent        CYGPKG_HAL_CORTEXM_KINETIS
    define_header hal_cortexm_kinetis_kwikstik.h
    include_dir   cyg/hal
    hardware

    requires      { is_active(CYGPKG_HAL_FREESCALE_EDMA) implies
        (CYGNUM_HAL_FREESCALE_EDMA_CHAN_NUM == 16) }

    requires      { CYGHWR_HAL_CORTEXM_KINETIS_SUBFAM == 40 }
    requires      { CYGHWR_HAL_CORTEXM_KINETIS_FPU == "D" }
    requires      { CYGHWR_HAL_CORTEXM_SYSTICK_CLK_SOURCE == "INTERNAL" }
    requires      { CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT_IS == "XTAL" ||
                    CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT_IS == "RTC" }
    requires      { CYGHWR_HAL_CORTEXM_KINETIS_FLEXNVM_DEFAULT == "X" }
    requires      { CYGHWR_HAL_CORTEXM_KINETIS_FLASH_NAME_DEFAULT == 256 }
    requires      { CYGHWR_HAL_CORTEXM_KINETIS_FLEXNVM == "X"
                    implies CYGHWR_HAL_KINETIS_FLEXRAM_SIZE == 4096 }

    implements    CYGINT_IO_SERIAL_FREESCALE_UART5
    implements    CYGINT_IO_FREESCALE_I2C1
    implements    CYGINT_HAL_FREESCALE_UART5
    implements    CYGINT_HAL_CORTEXM_KINETIS_RTC


    description   "
        The Freescale KwikStik Platform HAL package provides
        the support needed to run eCos on the KwikStik development
        system. This package can also be used for other boards that
        employ a controller from Kinetis families."

    compile       kwikstik_misc.c

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_cortexm_kinetis_kwikstik.h>"
        puts $::cdl_header "#define HAL_PLATFORM_CPU    \"Cortex-M4\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Freescale KwikStik\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
    }

    cdl_component CYG_HAL_STARTUP_ENV {
        display "Startup type"
        flavor data
        no_define
        calculated {
            !CYG_HAL_STARTUP_PLF ? CYG_HAL_STARTUP :
            ((CYG_HAL_STARTUP_PLF == "ByVariant") ?
            (CYG_HAL_STARTUP . "(Variant)") :
            (CYG_HAL_STARTUP . "(Platform)"))
        }
        description "
            Startup type configuration defines the system memory layout.
            Startup type  can be defined by the variant (CYG_HAL_STARTUP_VAR)
            or a platform (CYG_HAL_STARTUP_PLF). If CYG_HAL_STARTUP_PLF
            is defined and not equal to 'ByVariant' then it shall
            override CYG_HAL_STARTUP_VAR."
    }

    cdl_option CYGHWR_HAL_CORTEXM_KINETIS_PLF_XTAL_OR_OSC_FREQ {
        display "Platform Reference Clock Frequency"
        flavor data
        parent CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT
        active_if { CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT_IS == "OSC" ||
                   CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT_IS == "XTAL" }
        default_value 4000000
        legal_values { 32768 4000000 }
    }

    cdl_option CYGHWR_HAL_CORTEXM_KINETIS_PLF_OSC_CAP {
        display "Platform requred XTAL || C \[pF\]"
        flavor bool
        default_value { CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT_IS == "XTAL" }
        parent CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT
        active_if { CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT_IS == "XTAL" }
        requires { CYGHWR_HAL_CORTEXM_KINETIS_OSC_CAP == 0 }
    }

    cdl_option CYGHWR_HAL_CORTEXM_KINETIS_PLF_RTC {
        display "Platform requred RTC XTAL || C \[pF\]"
        flavor bool
        default_value 0
        parent CYGHWR_HAL_CORTEXM_KINETIS_RTC
        requires { CYGHWR_HAL_CORTEXM_KINETIS_RTC_OSC_CAP == 20 }
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        legal_values 0 to 2
        default_value   1
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The TWR board has one serial port fitted to RS232 connector.
            This optionchooses which port will be used to connect to a host
            running GDB."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
        display          "Diagnostic serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The TWR has one serial port fitted to RS232 connector.
            This option chooses which port will be used for diagnostic output."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Console serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 38400
        description   "
            This option controls the default baud rate used for the
            console connection.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 38400
        description   "
            This option controls the default baud rate used for the
            GDB connection.
            Note: this should match the value chosen for the console
            port if the console and GDB port are the same."
    }

    cdl_component CYGHWR_HAL_DEVS_IRQ_PRIO_SCHEME {
        display "Interrupt priority scheme"
        flavor none
        description "Consolidated interrupt priority scheme setting."
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        no_define
        parent  CYGPKG_NONE
        description   "
        Global build options including control over
        compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-eabi" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGBLD_GLOBAL_WARNFLAGS . "-mcpu=cortex-m3 -mthumb -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions" }
            description   "
            This option controls the global compiler flags which are used to
            compile all packages by default. Individual packages may define
            options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-mcpu=cortex-m3 -mthumb -Wl,--gc-sections -Wl,-static -Wl,-n -g -nostdlib" }
            description   "
            This option controls the global linker flags. Individual
            packages may define options which override these global flags."
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" || CYG_HAL_STARTUP == "JTAG" }
        requires      { CYGDBG_HAL_CRCTABLE_LOCATION == "ROM" }
        description   "
            Enable this option if this program is to be used as a
            ROM monitor, i.e. applications will be loaded into RAM on the
            board, and this ROM monitor may process exceptions or interrupts
            generated from the application. This enables features such as
            utilizing a separate interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
        display       "Work with a ROM monitor"
        flavor        booldata
        legal_values  { "Generic" "GDB_stubs" }
        default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "RAM" }
        description   "
            Support can be enabled for different varieties of ROM monitor.
            This support changes various eCos semantics such as the encoding
            of diagnostic output, or the overriding of hardware interrupt
            vectors.
            Firstly there is \"Generic\" support which prevents the HAL
            from overriding the hardware vectors that it does not use, to
            instead allow an installed ROM monitor to handle them. This is
            the most basic support which is likely to be common to most
            implementations of ROM monitor.
            \"GDB_stubs\" provides support when GDB stubs are included in
            the ROM monitor or boot ROM."
    }


    cdl_component CYGBLD_HAL_CORTEXM_KWIKSTIK_GDB_STUBS {
        display "Create StubROM SREC and binary files"
        active_if CYGBLD_BUILD_COMMON_GDB_STUBS
        no_define
        calculated 1
        requires { CYG_HAL_STARTUP == "ROM" }

        make -priority 325 {
            <PREFIX>/bin/stubrom.srec : <PREFIX>/bin/gdb_module.img
            $(OBJCOPY) -O srec $< $@
        }
        make -priority 325 {
            <PREFIX>/bin/stubrom.bin : <PREFIX>/bin/gdb_module.img
            $(OBJCOPY) -O binary $< $@
        }

        description "
            This component causes the ELF image generated by the
            build process to be converted to S-Record and binary
            files."
    }
}
