# ====================================================================
#
#      hal_h8300_h8s_sim.cdl
#
#      H8S SIM HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      ysato
# Original data:  bartv
# Contributors:
# Date:           2003-01-01
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_H8300_H8S_SIM {
    display  "H8S simulator"
    parent        CYGPKG_HAL_H8300
    requires CYGPKG_HAL_H8300_H8S
    implements CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    define_header hal_h8300_h8s_sim.h
    include_dir   cyg/hal
    description   "
           The minimal simulator HAL package is provided for use when
           only a simple simulation of the processor architecture is
           desired, as opposed to detailed simulation of any specific
           board. In particular it is not possible to simulate any of
           the I/O devices, so device drivers cannot be used."

    compile       hal_diag.c plf_misc.c delay_us.S

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H <pkgconf/hal_h8300_h8s.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_h8300_h8s_sim.h>"

        puts $::cdl_header "#define CYG_HAL_H8300"
	puts $::cdl_header "#define CYGNUM_HAL_H8300_SCI_PORTS 1"
	puts $::cdl_header "#define CYGHWR_HAL_VECTOR_TABLE 0xfff000"
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM"}
        default_value {"RAM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
            Only supports RAM startup."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   1
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           The CQ/7708 board has only one serial port. This option
           chooses which port will be used to connect to a host
           running GDB."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
	cdl_option CYGNUM_HAL_H8300_RTC_PRESCALE {
            display       "Real-time clock base prescale"
            flavor        data
	    calculated    8192
	}
        # Isn't a nice way to handle freq requirement!
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    10
        }
    }

    cdl_option CYGHWR_HAL_H8300_CPG_INPUT {
        display "OSC/Clock Freqency"
	flavor	data
	default_value 8000000
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "h8300-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGBLD_GLOBAL_WARNFLAGS . " -g -O2 -ms -mint32 -fsigned-char -fdata-sections -fno-rtti -fno-exceptions " }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-g -nostdlib -Wl,--gc-sections -Wl,-static -mrelax -ms -mint32" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { "h8300_h8s_sim_ram" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { "<pkgconf/mlt_h8300_h8s_sim_ram.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { "<pkgconf/mlt_h8300_h8s_sim_ram.h>" }
        }
    }
    cdl_option CYGHAL_PLF_SCI_BASE {
        display "SCI Base address"
        flavor data
	default_value 0xffff78
        description   "
            Used SCI Channel base address."
    }
}
