##==========================================================================
##
##      kinetis_irq_scheme.cdl
##
##      Cortex-M Freescale Kinetis IRQ configuration data
##
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2010, 2011 Free Software Foundation, Inc.                  
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##==========================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):    Ilija Kocho <ilijak@siva.com.mk>
## Date:         2010-12-05
##
######DESCRIPTIONEND####
##
##==========================================================================


#    cdl_component CYGHWR_HAL_DEVS_IRQ_PRIO_SCHEME_VAR {
#        display "Variant IRQ priority defaults"
#        no_define
#        flavor none
#        parent CYGHWR_HAL_DEVS_IRQ_PRIO_SCHEME
#        description "
#            Interrupt priorities defined by Kinetis variant"

        cdl_option CYGNUM_HAL_KERNEL_COUNTERS_CLOCK_ISR_DEFAULT_PRIORITY_SP {
            display       "Clock IRQ priority"
            flavor        data
            no_define
            default_value 0xE0
            description   "Set clock ISR priority. Default setting is lowest priority."
            legal_values { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80
                0x90 0xA0 0xB0 0xC0 0xD0 0xE0 }

        }

        cdl_option CYGNUM_DEVS_ETH_FREESCALE_ENET0_INTPRIO_SP {
            display "Ethernet IRQ priority"
            flavor data
            no_define
            active_if CYGPKG_DEVS_ETH_FREESCALE_ENET
            legal_values { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80
                0x90 0xA0 0xB0 0xC0 0xD0 0xE0 }
            default_value 0xE0
        }

        cdl_component CYGHWR_HAL_DEVS_IRQ_PRIO_SCHEME_UART {
            display "UART IRQ priorities"
            flavor none
            no_define

            cdl_option CYGNUM_IO_SERIAL_FREESCALE_UART0_INT_PRIORITY_SP {
                display "UART0 interrupt priority"
                flavor data
                no_define
                active_if CYGPKG_IO_SERIAL_FREESCALE_UART0
                legal_values { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80
                    0x90 0xA0 0xB0 0xC0 0xD0 0xE0 }
                default_value 0x80
            }

            cdl_option CYGNUM_IO_SERIAL_FREESCALE_UART1_INT_PRIORITY_SP {
                display "UART1 interrupt priority"
                flavor data
                no_define
                active_if CYGPKG_IO_SERIAL_FREESCALE_UART1
                legal_values { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80
                    0x90 0xA0 0xB0 0xC0 0xD0 0xE0 }
                default_value 0x80
            }

            cdl_option CYGNUM_IO_SERIAL_FREESCALE_UART2_INT_PRIORITY_SP {
                display "UART2 interrupt priority"
                flavor data
                no_define
                active_if CYGPKG_IO_SERIAL_FREESCALE_UART2
                legal_values { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80
                    0x90 0xA0 0xB0 0xC0 0xD0 0xE0 }
                default_value 0x80
            }

            cdl_option CYGNUM_IO_SERIAL_FREESCALE_UART3_INT_PRIORITY_SP {
                display "UART3 interrupt priority"
                flavor data
                no_define
                active_if CYGPKG_IO_SERIAL_FREESCALE_UART3
                legal_values { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80
                    0x90 0xA0 0xB0 0xC0 0xD0 0xE0 }
                default_value 0x80
            }

            cdl_option CYGNUM_IO_SERIAL_FREESCALE_UART4_INT_PRIORITY_SP {
                display "UART4 interrupt priority"
                flavor data
                no_define
                active_if CYGPKG_IO_SERIAL_FREESCALE_UART4
                legal_values { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80
                    0x90 0xA0 0xB0 0xC0 0xD0 0xE0 }
                default_value 0x80
            }

            cdl_option CYGNUM_IO_SERIAL_FREESCALE_UART5_INT_PRIORITY_SP {
                display "UART5 interrupt priority"
                flavor data
                no_define
                active_if CYGPKG_IO_SERIAL_FREESCALE_UART5
                legal_values { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80
                    0x90 0xA0 0xB0 0xC0 0xD0 0xE0 }
                default_value 0x80
            }
        }

        cdl_component CYGHWR_HAL_DEVS_IRQ_PRIO_SCHEME_DSPI {
            display "DSPI IRQ priorities"
            flavor none
            no_define

            cdl_option CYGNUM_DEVS_SPI_FREESCALE_DSPI0_ISR_PRI_SP {
                display "DSPI bus 0 interrupt priority"
                flavor data
                no_define
                active_if CYGHWR_DEVS_SPI_FREESCALE_DSPI0
                legal_values { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80
                    0x90 0xA0 0xB0 0xC0 0xD0 0xE0 }
                default_value 0xD0
            }

            cdl_option CYGNUM_DEVS_SPI_FREESCALE_DSPI1_ISR_PRI_SP {
                display "DSPI bus 1 interrupt priority"
                flavor data
                no_define
                active_if CYGHWR_DEVS_SPI_FREESCALE_DSPI1
                legal_values { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80
                    0x90 0xA0 0xB0 0xC0 0xD0 0xE0 }
                default_value 0xD0
            }

            cdl_option CYGNUM_DEVS_SPI_FREESCALE_DSPI2_ISR_PRI_SP {
                display "DSPI bus 2 interrupt priority"
                flavor data
                no_define
                active_if CYGHWR_DEVS_SPI_FREESCALE_DSPI2
                legal_values { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80
                    0x90 0xA0 0xB0 0xC0 0xD0 0xE0 }
                default_value 0xD0
            }
        }
        
        cdl_component CYGHWR_HAL_DEVS_IRQ_PRIO_SCHEME_I2C {
            display "I2C interrupt priorities"
            flavor none
            no_define
            
            for { set ::bus 0 } { $::bus < 2 } { incr ::bus } {
                
                cdl_option CYGNUM_DEVS_FREESCALE_I2C[set ::bus]_IRQ_PRIORITY {
                    display       "I2C bus [set ::bus] interrupt priority"
                    flavor        data
                    active_if     CYGHWR_DEVS_FREESCALE_I2C[set ::bus]
                    default_value 0x90
                    legal_values  { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80 
                        0x90  0xA0 0xB0 0xC0 0xD0 0xE0 }
                }
            }
        }

#    }


# EOF kinetis_irq_scheme.cdl
