#====================================================================
#
#      moab_eth_drivers.cdl
#
#      Hardware specifics for TAMS MOAB ethernet
#
#====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:   gthomas
# Date:           2003-08-19
#
#####DESCRIPTIONEND####
#
#====================================================================

cdl_package CYGPKG_DEVS_ETH_POWERPC_MOAB {
    display       "TAMS MOAB (PPC405GPr) ethernet support"
    description   "Hardware specifics for TAMS MOAB ethernet"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_HAL_POWERPC 
    active_if	  CYGPKG_HAL_POWERPC_PPC40x

    requires      CYGPKG_DEVS_ETH_POWERPC_PPC405
    requires      CYGHWR_DEVS_ETH_PHY_DP8384X
    requires      CYGPKG_HAL_POWERPC_MOAB

    # FIXME: This really belongs in the NS DP83816 package
    cdl_interface CYGINT_DEVS_ETH_NS_DP83816_REQUIRED {
        display   "NS DP83816 ethernet driver required"
    }

    cdl_component CYGHWR_DEVS_ETH_POWERPC_MOAB_ETH0 {
        display       "Include eth0 ethernet device"
        default_value 1
        description   "
          This option controls whether a driver for eth0
          is included in the resulting system."
        implements    CYGHWR_NET_DRIVERS
        implements    CYGHWR_NET_DRIVER_ETH0
        implements    CYGHWR_DEVS_ETH_POWERPC_PPC405_NET_DRIVERS
    }

    cdl_component CYGHWR_DEVS_ETH_POWERPC_MOAB_ETH1 {
        display       "Include eth1 ethernet device"
        default_value 1
        description   "
          This option controls whether a driver for eth1
          is included in the resulting system."
        implements    CYGHWR_NET_DRIVERS
        implements    CYGHWR_NET_DRIVER_ETH1
        requires      CYGHWR_DEVS_ETH_POWERPC_MOAB_ETH0

        implements CYGINT_DEVS_ETH_NS_DP83816_REQUIRED
	
        define_proc {
            puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
            puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_NS_DP83816_INL <cyg/io/moab_eth_dp83816.inl>"
            puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_NS_DP83816_CFG <pkgconf/devs_eth_powerpc_moab.h>"
            puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
        }

        cdl_option CYGNUM_DEVS_ETH_MOAB_DP83816_TxNUM {
            display       "Number of output buffers"
            flavor        data
            legal_values  2 to 64
            default_value 16
            description   "
                This option specifies the number of output buffer packets
                to be used for the NS DP83816 ethernet device."
        }
    
        cdl_option CYGNUM_DEVS_ETH_MOAB_DP83816_RxNUM {
            display       "Number of input buffers"
            flavor        data
            legal_values  2 to 64
            default_value 16
            description   "
                This option specifies the number of input buffer packets
                to be used for the NS DP83816 ethernet device."
        }
    }

    include_dir   cyg/io

    define_proc {
        puts $::cdl_system_header "#define CYGDAT_DEVS_PPC405_ETH_CDL <pkgconf/devs_eth_powerpc_moab.h>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_PPC405_ETH_INL <cyg/io/moab_eth.inl>"
    }
}
