# ====================================================================
#
#      microwindows.cdl
#
#      MicroWindows configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  jskov
# Contributors:
# Date:           2002-03-25
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_MICROWINDOWS {
    display       "MicroWindows"
    requires      CYGPKG_POSIX
    requires      CYGPKG_POSIX_TIMERS
    requires      CYGPKG_ISOINFRA
    requires      CYGINT_ISO_C_TIME_TYPES
    requires      CYGINT_ISO_STRERROR
    requires      CYGINT_ISO_ERRNO
    requires      CYGINT_ISO_ERRNO_CODES
    requires      CYGINT_ISO_MALLOC
    requires      CYGINT_ISO_STRING_BSD_FUNCS
    requires      CYGPKG_IO_FILEIO
    requires      CYGPKG_NET_STACK_INET
    description   "Microwindows."

    # Note: separating the stack implementation from the common support leads
    # to some rather incestious config file relationships.
    define_proc {
    }

    # FB drivers
    compile                                             \
        drivers/fblin16.c				\
        drivers/fblin1.c				\
        drivers/fblin24.c				\
        drivers/fblin2.c				\
        drivers/fblin32.c				\
        drivers/fblin4.c				\
        drivers/fblin8.c				\
        drivers/fb.c					\
        drivers/fbportrait_down.c			\
        drivers/fbportrait_left.c			\
        drivers/fbportrait_right.c			\
        drivers/genfont.c				\
        drivers/genmem.c

     # engine
     compile					\
        engine/devarc.c				\
        engine/devclip.c			\
        engine/devdraw.c			\
        engine/devfont.c			\
        engine/devimage.c			\
        engine/devkbd.c				\
        engine/devlist.c			\
        engine/devmouse.c			\
        engine/devopen.c			\
        engine/devpal1.c			\
        engine/devpal2.c			\
        engine/devpal4.c			\
        engine/devpal8.c			\
        engine/devpoly.c			\
        engine/devrgn2.c			\
        engine/devrgn.c				\
        engine/devtimer.c			\
        engine/error.c				\
        engine/selfont.c

     # NANO X
     compile					\
        nanox/srvmain.c				\
        nanox/srvfunc.c				\
        nanox/srvutil.c				\
        nanox/srvevent.c			\
        nanox/srvclip.c				\
        nanox/srvnet.c				\
        nanox/clientfb.c			\
        nanox/client.c				\
        nanox/error.c				\
        nanox/nxdraw.c				\
        nanox/nxproto.c				\
        nanox/nxutil.c

     # FONTS
     compile					\
        fonts/helvB10.c				\
        fonts/helvB12.c				\
        fonts/helvR10.c				\
        fonts/rom8x16.c				\
        fonts/rom8x8.c				\
        fonts/symbol.c				\
        fonts/winFreeSansSerif11x13.c		\
        fonts/winFreeSystem14x16.c		\
        fonts/X5x7.c				\
        fonts/X6x13.c

    # eCos stuff
    cdl_component CYGBLD_MICROWINDOWS_ECOS {
        display   "Build MicroWindows eCos support"
        default_value 0

        # These files are unique to eCos
        compile ecos/ecos_init.c 
        compile -library=libextras.a ecos/nanox_thread.c

        cdl_option CYGBLD_MICROWINDOWS_ECOS_APP {
            display  "Build complete eCos+MicroWindows application"
            default_value 0
            make -priority 320 {
                <PREFIX>/bin/ecos_mw.elf : $(PREFIX)/lib/target.ld $(PREFIX)/lib/vectors.o $(PREFIX)/lib/libtarget.a $(PREFIX)/lib/libextras.a $(REPOSITORY)/$(PACKAGE)/src/ecos/ecos_app.c
                        @sh -c "mkdir -p $(dir $@)"
                        $(CC) -c $(INCLUDE_PATH) $(CFLAGS) -o $(PREFIX)/lib/ecos_app.o $(REPOSITORY)/$(PACKAGE)/src/ecos/ecos_app.c
                        $(CC) $(LDFLAGS) -L$(PREFIX)/lib -Ttarget.ld -o $@ $(PREFIX)/lib/ecos_app.o
            }
            
        }
    }

    # eCos VNC server drivers
    cdl_option CYGBLD_MICROWINDOWS_VNC_DRIVERS {
        display   "Build MicroWindows VNC server drivers"
        default_value 0
        description \
            "This option builds the drivers for the VNC server.  The VNC server
             then provides a virtual screen, keyboard and mouse for MicroWindows."

        compile                     \
            drivers/scr_vnc_ecos.c  \
            drivers/kbd_vnc_ecos.c  \
            drivers/mou_vnc_ecos.c
            
        requires CYGBLD_MICROWINDOWS_ECOS
        requires CYGBLD_MICROWINDOWS_NANOWM
        requires CYGPKG_VNC_SERVER
        requires !CYGBLD_MICROWINDOWS_ARM_DRIVERS
        requires CYGPKG_VNC_SERVER_BUILD_MOUSE_DRIVER
        requires CYGPKG_VNC_SERVER_BUILD_KEYBOARD_DRIVER
    }

    # eCos ARM drivers
    cdl_option CYGBLD_MICROWINDOWS_ARM_DRIVERS {
        display   "Build MicroWindows ARM drivers"
        default_value CYGPKG_HAL_ARM

        compile					\
            drivers/scr_ecos.c                  \
            drivers/kbd_ipaq.c			\
            drivers/mou_ipaq.c


        requires CYGBLD_MICROWINDOWS_ECOS
        requires CYGBLD_MICROWINDOWS_NANOWM
        requires CYGBLD_MICROWINDOWS_NXKBD
        requires CYGBLD_MICROWINDOWS_NANOX_DEMOS

        # This should come from the HAL
        requires { !CYGPKG_HAL_ARM_SA11X0_IPAQ || is_substr(CYGPKG_MICROWINDOWS_CFLAGS_ADD, " -DMWPIXEL_FORMAT=MWPF_TRUECOLOR565") }
        requires { !CYGPKG_HAL_ARM_ARM9_AAED2000 || is_substr(CYGPKG_MICROWINDOWS_CFLAGS_ADD, " -DMWPIXEL_FORMAT=MWPF_TRUECOLOR555") }

    }

    cdl_component CYGPKG_MICROWINDOWS_PC {
	display     "Build options for PC hardware"
	flavor      none
    active_if   (CYGPKG_HAL_I386_PCMB && !CYGBLD_MICROWINDOWS_VNC_DRIVERS)
	compile     drivers/ps2kbdmou_ecos.c
	
	requires CYGBLD_MICROWINDOWS_ECOS
	
	cdl_option CYGIMP_MICROWINDOWS_PCSVGA32 {
	    display "Assume 32 bits per pixel, RGB == 0888"
	    description \
		"This mode can be used when building for a standard PC,
	         where bootstrap is handled via RedBoot. A custom version
	         of RedBoot is required, configured to switch the graphics
	         card to a suitable resolution before the processor enters
	         protected mode. A VESA-compliant video BIOS is used for
	         this. The graphics mode should be 32 bits per pixel true-color."

	    implements CYGINT_MICROWINDOWS_PC_DRIVER
	    default_value 1
	    compile drivers/scr_ecospcsvga.c
	    requires { is_substr(CYGPKG_MICROWINDOWS_CFLAGS_ADD, " -DMWPIXEL_FORMAT=MWPF_TRUECOLOR0888 ") }
	    requires { !is_substr(CYGPKG_MICROWINDOWS_CFLAGS_ADD, " -DMWPIXEL_FORMAT=MWPF_TRUECOLOR565 ") }
	    requires { !is_substr(CYGPKG_MICROWINDOWS_CFLAGS_ADD, " -DMWPIXEL_FORMAT=MWPF_PALETTE ") }
	}
	
	cdl_option CYGIMP_MICROWINDOWS_PCSVGA16 {
	    display "Assume 16 bits per pixel, RGB == 565"
	    description \
		"This mode can be used when building for a standard PC,
	         where bootstrap is handled via RedBoot. A custom version
	         of RedBoot is required, configured to switch the graphics
	         card to a suitable resolution before the processor enters
	         protected mode. A VESA-compliant video BIOS is used for
	         this. The graphics mode should be 16 bits per pixel true-color."

	    implements CYGINT_MICROWINDOWS_PC_DRIVER
	    default_value 0
	    compile drivers/scr_ecospcsvga.c
	    requires { !is_substr(CYGPKG_MICROWINDOWS_CFLAGS_ADD, " -DMWPIXEL_FORMAT=MWPF_TRUECOLOR0888 ") }
	    requires { is_substr(CYGPKG_MICROWINDOWS_CFLAGS_ADD, " -DMWPIXEL_FORMAT=MWPF_TRUECOLOR565 ") }
	    requires { !is_substr(CYGPKG_MICROWINDOWS_CFLAGS_ADD, " -DMWPIXEL_FORMAT=MWPF_PALETTE ") }
	}
	
	cdl_option CYGIMP_MICROWINDOWS_PCVGA {
	    display "Build for VGA hardware"
	    description \
		"This driver manipulates VGA hardware directly, rather than
	         going via the video BIOS. Only a limited resolution of
	         640x480 with 4 bits per pixel is available. The driver
	         does not implement all required microwindows functionality."

	    implements CYGINT_MICROWINDOWS_PC_DRIVER
	    default_value 0
	    compile drivers/scr_bios.c drivers/vgainit.c drivers/vgaplan4.c drivers/memplan4.c
	    requires { is_substr(CYGPKG_MICROWINDOWS_CFLAGS_ADD, " -DMWPIXEL_FORMAT=MWPF_PALETTE ") }
	    requires { !is_substr(CYGPKG_MICROWINDOWS_CFLAGS_ADD, " -DMWPIXEL_FORMAT=MWPF_TRUECOLOR0888 ") }
	}
	
	cdl_interface CYGINT_MICROWINDOWS_PC_DRIVER {
	    display "Number of active PC graphics drivers"
	    requires { CYGINT_MICROWINDOWS_PC_DRIVER == 1 }
	}
    }
    

    # Nano WM
    cdl_option CYGBLD_MICROWINDOWS_NANOWM {
        display   "Build MicroWindows NANOWM"
        default_value 0

        compile					\
            demos/nanowm/nanowm.c			\
            demos/nanowm/events.c			\
            demos/nanowm/wlist.c			\
            demos/nanowm/clients.c			\
            demos/nanowm/actions.c                      
        compile -library=libextras.a ecos/nanowm_thread.c
    }

    # keyboard
    cdl_option CYGBLD_MICROWINDOWS_NXKBD {
        display   "Build MicroWindows NXKBD"
        default_value 0

        compile					\
            demos/nxkbd/nxkbd.c			\
            demos/nxkbd/srvconn.c			\
            demos/nxkbd/keynorm.c			\
            demos/nxkbd/keyctrl.c			\
            demos/nxkbd/keyshft.c			\
            demos/nxkbd/keynum.c
    }

    # keyboard
    cdl_component CYGBLD_MICROWINDOWS_NANOX_DEMOS {
        display   "Build MicroWindows NanoX demos"
        default_value 0

        cdl_option CYGBLD_MICROWINDOWS_NANOX_DEMOS_WORLD {
            display "Include 'world' demo"
            default_value 0
            no_define
            compile demos/nanox/world.c 
            compile -library=libextras.a ecos/world_thread.c
        }

        cdl_option CYGBLD_MICROWINDOWS_NANOX_DEMOS_NTETRIS {
            display "Include 'nano-tetris' demo"
            default_value 0
            no_define
            compile demos/nanox/ntetris.c 
            compile -library=libextras.a ecos/ntetris_thread.c
        }
    }

    cdl_component CYGPKG_MICROWINDOWS_OPTIONS {
        display "Build options"
        flavor  none
        no_define
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_MICROWINDOWS_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-I$(PREFIX)/include/microwin -D__ECOS=1 -DMSDOS=0 -DELKS=0 -D__rtems__=0 -D_MINIX=0 -DNOTYET=0 -DUNIX=1 -DHAVE_FILEIO -DHAVE_BMP_SUPPORT=1 -DHAVE_PNM_SUPPORT=1 -DHAVE_XPM_SUPPORT=1 -DxHAVE_JPEG_SUPPORT=1 -DHAVESELECT=1" }
            description   "
                This option modifies the set of compiler flags for
                building the MicroWindows package.
                These flags are used in addition to the set of global flags."
        }

        cdl_option CYGPKG_MICROWINDOWS_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the MicroWindows package.
                These flags are removed from the set of global flags
                if present."
        }
    }
}
