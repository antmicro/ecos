#==========================================================================
# 
#       i2c_xc7z.cdl
# 
#       eCos configuration data for the Xilinx Zynq i2c device
# 
#==========================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
#==========================================================================
######DESCRIPTIONBEGIN####
# 
# Author(s):    Ant Micro <www.antmicro.com>
# Date:         2012-07-23
# Purpose:      
# Description:  I2C configuration data for Xilinx Zynq
# 
#####DESCRIPTIONEND####
# 
#==========================================================================


cdl_package CYGPKG_DEVS_I2C_ARM_XC7Z {
    display       "Xilinx Zynq I2C driver"

    parent        CYGPKG_IO_I2C
    active_if     CYGPKG_IO_I2C
    
    implements    CYGINT_I2C_HW_IMPLEMENTATIONS
    implements    CYGINT_I2C_RESETS_ON_TIMEOUT

    description   "
        Xilinx Zynq I2C driver"

    compile       i2c_xc7z.c     
    include_dir   cyg/io

    cdl_option CYGPKG_DEVS_I2C_ARM_XC7Z_INTERFACE {
        display "Used I2C interface"
        flavor data
        default_value 1
        legal_values {0 1}
	    description "
		This option defines which hardware I2C interface
		(0 or 1) will be used."
    }
   
    cdl_option CYGPKG_DEVS_I2C_ARM_XC7Z_PCLK {
        display "CPU input clock in Hz"
        flavor data
        default_value { 111000000 }
	    description "
		Value of the CPU input clock in Hz.
		It is not I2C SCL frequency!"
    }
    
    cdl_option CYGBLD_DEVS_I2C_ARM_XC7Z_STD_TEST {
        display       "Build Zynq I2C test"
        flavor        bool
        no_define
        default_value 0
        description   "
            This option enables the building of the Xilinx Zynq I2C test."
    }

    cdl_option CYGPKG_DEVS_I2C_ARM_XC7Z_TESTS {
        display         "I2C standard test"
        flavor          data
        no_define
        calculated      { CYGBLD_DEVS_I2C_ARM_XC7Z_STD_TEST ? "tests/i2ctest" : "" } 
    }
}



