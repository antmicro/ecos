# ====================================================================
#
#      spi_xc7z.cdl
#
#      Xilinx XC7Z020 (ARM) SPI driver configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2009 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):    Antmicro Ltd <www.antmicro.com>, Artur Łącki <alacki93@gmail.com>
# Date:         2015-08-31
# Purpose:
# Description:    SPI configuration data for Xilinx Zynq
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_SPI_ARM_XC7Z {
    parent        CYGPKG_IO_SPI
    active_if     CYGPKG_IO_SPI
    display       "Xilinx Zynq SPI driver"
    requires      CYGPKG_HAL_ARM_XC7Z020
    requires      CYGPKG_HAL_ARM
    requires      CYGPKG_ERROR
    hardware
    include_dir   cyg/io
    compile       spi_xc7z.c
    compile       -library=libextras.a spi_xc7z_init.cxx

    cdl_option CYGHWR_DEVS_SPI_ARM_XC7Z_BUS0 {
        display       "Enable support for SPI bus 0"
        flavor        bool
        default_value 1
    }

    cdl_option CYGHWR_DEVS_SPI_ARM_XC7Z_BUS1 {
        display       "Enable support for SPI bus 1"
        flavor        bool
        default_value 1
    }
}


# EOF spi_xc7z.cdl
