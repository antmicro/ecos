# ====================================================================
#
#      i2c_mcf52xx.cdl
#
#      eCos MCF52xx I2C configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2005, 2006 Free Software Foundation, Inc.                  
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Uwe Kindler
# Contributors:   Bart Veer
# Date:           2005-10-23
#
#####DESCRIPTIONEND####
# ====================================================================


cdl_package CYGPKG_DEVS_I2C_MCF52xx {
    display         "I2C driver for coldfire MCF52xx family"
    doc             ref/devs-i2c-m68k-mcf52xx-part.html

    parent          CYGPKG_IO_I2C
    active_if       CYGPKG_IO_I2C
    active_if       CYGPKG_HAL_M68K_MCF52xx

    description   "
           This package provides a generic I2C device driver for the on-chip
           I2C modules in MCF52xx ColdFire processors."

    include_dir     cyg/io
    compile 	    i2c_mcf52xx.c

    cdl_option CYGHWR_DEVS_I2C_MCF52xx_MULTIPLE_BUSES {
	display		"Target hardware may have multiple MCF52xx I2C buses"
	flavor		bool
	default_value	0
	description "
            The MCF52xx I2C driver can support multiple I2C bus devices, but
          typically the coldfire processor only provides a single device. By
          default the driver assumes only a single device is present and will
          optimize for that case, using constant definitions provided by the
          platform HAL rather than per-device structure fields. If the hardware
          has multiple I2C bus devices, or if a singleton bus is instantiated
          by some other package and hence the platform HAL cannot provide the
          necessary definitions, then this option should be enabled."
    }
    
    cdl_component CYGPKG_DEVS_I2C_MCF52xx_OPTIONS {
        display 	"I2C driver build options"
        flavor  	none
	active_if	{ CYGINT_DEVS_I2C_MCF52xx_BUS_DEVICES > 0 }
        description   "
	    Package specific build options including control over
	    compiler flags used only in building the MCF52xx I2C
            bus driver."

        cdl_option CYGPKG_DEVS_I2C_MCF52xx_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the MCF52xx I2C bus driver. These flags are
                used in addition to the set of global flags."
        }

        cdl_option CYGPKG_DEVS_I2C_MCF52xx_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the MCF52xx I2C bus driver. These flags are
                removed from the set of global flags if present."
        }
    }
}
