# ====================================================================
#
#      ser_sh_se77x9.cdl
#
#      eCos serial SH/SE77X9 configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:
# Date:           2001-06-18
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_SH_SE77X9 {
    display       "SH3 SE77X9 serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_SH_SH77X9_SE77X9

    requires      CYGPKG_ERROR
    include_dir   cyg/io

    description   "
        This option enables the serial device drivers for the
        Hitachi SH3 SE77X9 board, based on the generic SH SCI driver."


    # FIXME: This really belongs in the SH_SCIF package
    cdl_interface CYGINT_IO_SERIAL_SH_SCIF_REQUIRED {
        display   "SH SCI driver required"
    }

    # FIXME: This really belongs in the GENERIC_16X5X package
    cdl_interface CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED {
        display   "Generic 16x5x serial driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_INL <cyg/io/sh_sh3_se77x9_16x5x.inl>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_CFG <pkgconf/io_serial_sh_se77x9.h>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_SH_SCIF_INL <cyg/io/sh_sh3_se77x9_scif.inl>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_SH_SCIF_CFG <pkgconf/io_serial_sh_se77x9.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

    cdl_component CYGPKG_IO_SERIAL_SH_SE77X9_COM1 {
        display       "SH SE77X9 serial 1 driver (SuperIO)"
        flavor        bool
        calculated    0
        description   "
            This option includes the serial device driver for the COM1
            port. FIXME: Disabled due to being broken."

        implements CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED
        implements CYGINT_IO_SERIAL_FLOW_CONTROL_HW
        implements CYGINT_IO_SERIAL_LINE_STATUS_HW

        cdl_option CYGDAT_IO_SERIAL_SH_SE77X9_COM1_NAME {
            display       "Device name for COM1"
            flavor        data
            default_value {"\"/dev/ser1\""}
            description   "
                This option specifies the device name for COM1."
        }

        cdl_option CYGNUM_IO_SERIAL_SH_SE77X9_COM1_BAUD {
            display       "Baud rate for COM1"
            flavor        data
            legal_values  { 4800 9600 14400 19200 38400 57600 115200 }
            default_value 38400
            description   "
                This option specifies the default baud rate (speed)
                for the COM1 port."
        }

        cdl_option CYGNUM_IO_SERIAL_SH_SE77X9_COM1_BUFSIZE {
            display       "Buffer size for COM1"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers
                used for the COM1 port."
        }
    }

    # SCIF port
    cdl_component CYGPKG_IO_SERIAL_SH_SE77X9_COM2 {
        display       "SE77X9 serial, SCIF port 2 driver"
        flavor        bool
        default_value 1
        description   "
            This option includes the serial device driver for SCIF
            port 2."

        implements CYGINT_IO_SERIAL_SH_SCIF_REQUIRED
        implements CYGINT_IO_SERIAL_FLOW_CONTROL_HW
        implements CYGINT_IO_SERIAL_LINE_STATUS_HW

        cdl_option CYGDAT_IO_SERIAL_SH_SE77X9_COM2_NAME {
            display       "Device name"
            flavor        data
            default_value {"\"/dev/ser2\""}
            description   "
                This option specifies the device name for the serial
                port."
        }

        cdl_option CYGNUM_IO_SERIAL_SH_SE77X9_COM2_BAUD {
            display       "Baud rate"
            flavor        data
            legal_values  { 4800 9600 14400 19200 38400 57600 115200 }
            default_value 38400
            description   "
                This option specifies the default baud rate (speed)
                for the serial driver."
        }

        cdl_option CYGNUM_IO_SERIAL_SH_SE77X9_COM2_BUFSIZE {
            display       "Buffer size"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers
                used for the serial driver."
        }

        cdl_option CYGSEM_IO_SERIAL_SH_SE77X9_COM2_DMA {
            display       "Enable SCIF serial driver DMA"
            active_if     CYGINT_HAL_SH_DMA_CHANNELS
            implements    CYGINT_HAL_SH_DMA_CHANNELS_USED
            implements    CYGINT_IO_SERIAL_SH_SCIF_DMA
            default_value 1
            description   "
                Enable DMA for this port."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_SH_SE77X9_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        no_define
        active_if  CYGPKG_IO_SERIAL_SH_SE77X9_COM2

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"sh-se77x9\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_SER_DEV  CYGDAT_IO_SERIAL_SH_SE77X9_COM2_NAME"
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty2\""
        }
    }
}
# EOF ser_sh_se77x9.cdl
