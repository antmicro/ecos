##=============================================================================
##
##      spi_a2fxxx.cdl
##
##      Smartfusion Cortex-M3 SPI driver configuration options.
##
##=============================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008, 2009, 2011 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##=============================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):   ccoutand, updated for Smartfusion Cortex-M3
## Original(s): Chris Holgate
## Date:        2011-04-25
## Purpose:     Configure Smartfusion Cortex-M3 SPI driver.
##
######DESCRIPTIONEND####
##
##=============================================================================

cdl_package CYGPKG_DEVS_SPI_CORTEXM_A2FXXX {
    display       "Actel Smartfusion SPI driver"
    description   "
        This package provides SPI driver support for the Smartfusion Cortex-M3
        series of microcontrollers.
    "
    parent        CYGPKG_IO_SPI
    active_if     CYGPKG_IO_SPI
    requires      CYGPKG_HAL_CORTEXM_A2FXXX
    hardware
    include_dir   cyg/io
    compile       -library=libextras.a spi_a2fxxx.c

    cdl_option CYGDBG_DEVS_SPI_CORTEXM_A2FXXX_TRACE {
        display       "Display status messages during SPI operations"
        flavor        bool
        default_value 0
        description   "
           Selecting this option will cause the SPI driver to print status
           messages as various SPI operations are undertaken."
    }

    cdl_component CYGHWR_DEVS_SPI_CORTEXM_A2FXXX_BUS1 {
        display       "Actel Smartfusion SPI bus 1"
        description   "
            Enable SPI bus 1 on the A2FXXX device.
            "
        flavor        bool
        default_value false

        cdl_option CYGNUM_DEVS_SPI_CORTEXM_A2FXXX_BUS1_TX_DMA {
            display       "Transmit DMA channel number"
            flavor        data
            default_value 0
        }

        cdl_option CYGNUM_DEVS_SPI_CORTEXM_A2FXXX_BUS1_RX_DMA {
            display       "Receive DMA channel number"
            flavor        data
            default_value 1
        }

        cdl_option CYGDAT_DEVS_SPI_CORTEXM_A2FXXX_BUS1_TX_DMA_PRI {
            display       "Transmit DMA channel priority"
            legal_values  { "HIGH" "LOW" }
            flavor        data
            default_value { "HIGH" }
        }

        cdl_option CYGDAT_DEVS_SPI_CORTEXM_A2FXXX_BUS1_RX_DMA_PRI {
            display       "Receive DMA channel priority"
            legal_values  { "HIGH" "LOW" }
            flavor        data
            default_value { "HIGH" }
        }
    }

    cdl_component CYGHWR_DEVS_SPI_CORTEXM_A2FXXX_BUS2 {
        display       "Actel Smartfusion SPI bus 2"
        description   "
            Enable SPI bus 2 on the A2FXXX device.
        "
        flavor        bool
        default_value false

        cdl_option CYGNUM_DEVS_SPI_CORTEXM_A2FXXX_BUS2_TX_DMA {
            display       "Transmit DMA channel number"
            flavor        data
            default_value 2
        }

        cdl_option CYGNUM_DEVS_SPI_CORTEXM_A2FXXX_BUS2_RX_DMA {
            display       "Receive DMA channel number"
            flavor        data
            default_value 3
        }

        cdl_option CYGDAT_DEVS_SPI_CORTEXM_A2FXXX_BUS2_TX_DMA_PRI {
            display       "Transmit DMA channel priority"
            legal_values  { "HIGH" "LOW" }
            flavor        data
            default_value { "HIGH" }
        }

        cdl_option CYGDAT_DEVS_SPI_CORTEXM_A2FXXX_BUS2_RX_DMA_PRI {
            display       "Receive DMA channel priority"
            legal_values  { "HIGH" "LOW" }
            flavor        data
            default_value { "HIGH" }
        }
    }

    cdl_component CYGPKG_DEVS_SPI_CORTEXM_A2FXXX_OPTIONS {
        display "Actel Smartfusion SPI driver build options"
        flavor  none
        description   "
        Package specific build options including control over
        compiler flags used only in building this package,
        and details of which tests are built."

        cdl_option CYGPKG_DEVS_SPI_CORTEXM_A2FXXX_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the A2FXXX SPI driver. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_DEVS_SPI_CORTEXM_A2FXXX_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the A2FXXX SPI driver. These flags are removed from
                the set of global flags if present."
        }
    }

}
# EOF spi_a2fxxx.cdl
