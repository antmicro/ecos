# ====================================================================
#
#      hal_h8300_h8300h_sim.cdl
#
#      AKI3068NET board HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      yoshinori sato
# Original data:  bartv
# Contributors:   yoshinori sato
# Date:           2002-04-10
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_H8300_H8300H_AKI3068NET {
    display  "AKI3068NET"
    parent        CYGPKG_HAL_H8300
    requires CYGPKG_HAL_H8300_H8300H
    implements CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    define_header hal_h8300_h8300h_aki3068net.h
    include_dir   cyg/hal
    description   "
           The aki HAL package provides the support needed to run
           eCos on a Akizuki H8/3068 Network micom board." 

    compile       hal_diag.c plf_misc.c delay_us.S plf_ide.c

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H <pkgconf/hal_h8300_h8300h.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_h8300_h8300h_aki3068net.h>"
	puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_IO_H <cyg/hal/plf_io.h>"

        puts $::cdl_header "#define CYG_HAL_H8300"
	puts $::cdl_header "#define CYGNUM_HAL_H8300_SCI_PORTS 1"
	puts $::cdl_header "#define CYGHWR_HAL_VECTOR_TABLE 0xfffe20"
        puts $::cdl_header "#define HAL_PLATFORM_CPU    \"H8/300H\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Akizuki H8/3068 Network micom\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"ROM" "RAM"}
        default_value {"ROM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
           When targetting the AKI3068NET board it is possible to
           build the system for either RAM bootstrap or ROM bootstrap.
           RAM bootstrap generally requires that the board
           is equipped with ROMs containing a suitable ROM monitor or
           equivalent software that allows GDB to download the eCos
           application and extend Memory on to the board. 
           The ROM bootstrap typically
           requires that the eCos application be blown into EPROMs or
           equivalent technology."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   1
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           The AKI3068NET board has only one serial port. This option
           chooses which port will be used to connect to a host
           running GDB."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
        display          "Diagnostic serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           The CQ/7708 board has only one serial port.  This option
           chooses which port will be used for diagnostic output."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            default_value 1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
        }
	cdl_option CYGNUM_HAL_H8300_RTC_PRESCALE {
            display       "Real-time clock base prescale"
            flavor        data
	    calculated    8192
	}
        # Isn't a nice way to handle freq requirement!
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            default_value 10
        }
    }

    cdl_option CYGHWR_HAL_H8300_CPG_INPUT {
        display "OSC/Clock Freqency"
	flavor	data
	default_value 20000000
    }

    cdl_option CYGHWR_HAL_AKI3068NET_EXTRAM {
	display "Extend DRAM Using"
	flavor	bool
	default_value 1
    }

    cdl_option CYGHWR_HAL_AKI3068NET_IDE {
	display "IDE I/F expand"
	flavor	bool
	default_value 0
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "h8300-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGBLD_GLOBAL_WARNFLAGS . " -g -O2 -mh -mint32 -fsigned-char -fdata-sections -fno-rtti -fno-exceptions " }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-g -nostdlib -Wl,--gc-sections -Wl,-static -mrelax -mh -mint32" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "h8300_h8300h_aki3068net_ram" : \
                                                "h8300_h8300h_aki3068net_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_h8300_h8300h_aki3068net_ram.ldi>" : \
                                                    "<pkgconf/mlt_h8300_h8300h_aki3068net_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_h8300_h8300h_aki3068net_ram.h>" : \
                                                    "<pkgconf/mlt_h8300_h8300h_aki3068net_rom.h>" }
        }
    }

    cdl_component CYGHWR_AKI3068NET_IDE_OPTIONS {
        display "IDE Expand Setting"
        flavor  none
        parent  CYGPKG_NONE
	active_if CYGHWR_HAL_AKI3068NET_IDE
	implements CYGINT_HAL_PLF_IF_IDE
        description   "
	    IDE Expand Hardware Setting."

	cdl_option CYGHWR_HAL_IDE_REGISTER {
	    display "IDE Register base address"
	    flavor  data
	    default_value 0x600000
        }

        cdl_option CYGHWR_HAL_IDE_ALT_REGS {
	    display "IDE AlternateRegister base address"
	    flavor  data
	    default_value 0x600020
        }

        cdl_option CYGHWR_HAL_IDE_BUSWIDTH {
	    display "IDE bus width"
	    flavor  data
	    legal_values  {8 16}
	    default_value 8
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }
    cdl_option CYGHWR_HAL_H8300_VECTOR_ADDRESS {
        display       "Hook Vector Address"
        flavor        data
        default_value 0xfffd20
	active_if CYGSEM_HAL_H8300_VECTOR_HOOK
        parent        CYGPKG_HAL_ROM_MONITOR
        description   "
            Hooking Vector Table Address"
    }
    cdl_option CYGHAL_PLF_SCI_BASE {
        display "SCI Base address"
        flavor data
	default_value 0xffffb8
        description   "
            Used SCI Channel base address."
    }
    cdl_option CYGDAT_REDBOOT_H8300_LINUX_COMMAND_START {
        display        "Default kernel command line start address"
        flavor         data
        default_value  0x5ffe00
        description    "
           This option uClinux kernel command line start address of default."
    }

    cdl_option CYGDAT_REDBOOT_H8300_LINUX_BOOT_COMMAND_LINE {
        display        "Default command line"
        flavor         data
        default_value  { "console=/dev/ttySC1" }
        description    "
           This option uClinux kernel startup command line of default."
    }
}
