# ====================================================================
#
#      hal_arm.cdl
#
#      ARM architectural HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2014 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      bartv
# Original data:  gthomas
# Contributors:   jld
# Date:           1999-06-13
#
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_HAL_ARM {
    display       "ARM architecture"
    parent        CYGPKG_HAL
    hardware
    include_dir   cyg/hal
    define_header hal_arm.h
    description   "
        The ARM architecture HAL package provides generic
        support for this processor architecture. It is also
        necessary to select a specific target platform HAL
        package."

    implements    CYGINT_PROFILE_HAL_MCOUNT

    compile       hal_misc.c context.S arm_stub.c hal_syscall.c

    # The "-o file" is a workaround for CR100958 - without it the
    # output file would end up in the source directory under CygWin.
    # n.b. grep does not behave itself under win32
    make -priority 1 {
        arm.inc : <PACKAGE>/src/hal_mk_defs.c
        $(CC) $(ACTUAL_CFLAGS) $(INCLUDE_PATH) -Wp,-MD,arm.tmp -o hal_mk_defs.tmp -S $<
        fgrep .equ hal_mk_defs.tmp | sed s/#// > $@
        @echo $@ ": \\" > $(notdir $@).deps
        @tail -n +2 arm.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm arm.tmp hal_mk_defs.tmp
    }

    make {
        <PREFIX>/lib/vectors.o : <PACKAGE>/src/vectors.S
        $(CC) -Wp,-MD,vectors.tmp $(INCLUDE_PATH) $(ACTUAL_CFLAGS) -c -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail -n +2 vectors.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm vectors.tmp
    }

    make {
        <PREFIX>/lib/target.ld: <PACKAGE>/src/arm.ld
        $(CC) -E -P -Wp,-MD,target.tmp -xc $(INCLUDE_PATH) $(ACTUAL_CFLAGS) -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail -n +2 target.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm target.tmp
    }

    cdl_component CYGPKG_HAL_SMP_SUPPORT {
      display       "SMP support"
      default_value 0
      requires { CYGPKG_HAL_ARM_MARS_ZX3 != 0 }

      cdl_option CYGPKG_HAL_SMP_CPU_MAX {
          display       "Max number of CPUs supported"
          flavor        data
          active_if     { CYGPKG_HAL_SMP_SUPPORT == 1 }
          legal_values  2
          default_value 2
      }
    }

    cdl_interface CYGINT_HAL_ARM_THUMB_ARCH {
        display "The CPU architecture supports THUMB mode"
    }

    cdl_option CYGHWR_THUMB {
        display          "Enable Thumb instruction set"
        active_if        { CYGINT_HAL_ARM_THUMB_ARCH != 0 }
        default_value    0
        description      "
            Enable use of the Thumb instruction set."
    }

    # Note that when building a ROM monitor we include Thumb
    # interworking in order to support Thumb applications running
    # under a ARM ROM monitor.
    cdl_option CYGBLD_ARM_ENABLE_THUMB_INTERWORK {
        display       "Enable Thumb interworking compiler option"
        active_if        { CYGINT_HAL_ARM_THUMB_ARCH != 0 }
        default_value { (CYGHWR_THUMB || CYGSEM_HAL_ROM_MONITOR) }
        description "
            This option controls the use of -mthumb-interwork in the
            compiler flags. It defaults enabled in Thumb or ROM monitor
            configurations, but can be overridden for reduced memory
            footprint where interworking is not a requirement."
    }

    cdl_interface CYGINT_HAL_ARM_BIGENDIAN {
        display "The platform and architecture supports Big Endian operation"
    }

    cdl_option CYGHWR_HAL_ARM_BIGENDIAN {
        display          "Use big-endian mode"
        active_if        { CYGINT_HAL_ARM_BIGENDIAN != 0 }
        default_value    0
        description      "
            Use the CPU in big-endian mode."
    }

    cdl_option CYGBLD_ARCH_CFLAGS {
        display     "Architecture-specific compiler flags"
        parent      CYGBLD_GLOBAL_OPTIONS
        flavor      data
        no_define
        calculated  { (CYGHWR_THUMB ? " -mthumb " : "") .
            (CYGBLD_ARM_ENABLE_THUMB_INTERWORK ? " -mthumb-interwork " : " -mno-thumb-interwork ") .
            (CYGHWR_HAL_ARM_BIGENDIAN ? " -mbig-endian " : "")
        }
        requires    {  CYGHWR_THUMB &&  CYGBLD_ARM_ENABLE_THUMB_INTERWORK implies  is_substr(CYGBLD_GLOBAL_CFLAGS, " -mthumb ") &&
                                                                                   is_substr(CYGBLD_GLOBAL_CFLAGS, " -mthumb-interwork ") &&
                                                                                  !is_substr(CYGBLD_GLOBAL_CFLAGS, " -mno-thumb-interwork ") }
        requires    { !CYGHWR_THUMB &&  CYGBLD_ARM_ENABLE_THUMB_INTERWORK implies !is_substr(CYGBLD_GLOBAL_CFLAGS, " -mthumb ") &&
                                                                                   is_substr(CYGBLD_GLOBAL_CFLAGS, " -mthumb-interwork ") &&
                                                                                  !is_substr(CYGBLD_GLOBAL_CFLAGS, " -mno-thumb-interwork ") }
        requires    {  CYGHWR_THUMB && !CYGBLD_ARM_ENABLE_THUMB_INTERWORK implies  is_substr(CYGBLD_GLOBAL_CFLAGS, " -mthumb ") &&
                                                                                  !is_substr(CYGBLD_GLOBAL_CFLAGS, " -mthumb-interwork ") &&
                                                                                   is_substr(CYGBLD_GLOBAL_CFLAGS, " -mno-thumb-interwork ") }
        requires    { !CYGHWR_THUMB && !CYGBLD_ARM_ENABLE_THUMB_INTERWORK implies !is_substr(CYGBLD_GLOBAL_CFLAGS, " -mthumb ") &&
                                                                                  !is_substr(CYGBLD_GLOBAL_CFLAGS, " -mthumb-interwork ") &&
                                                                                   is_substr(CYGBLD_GLOBAL_CFLAGS, " -mno-thumb-interwork ") }
        requires    {  CYGHWR_HAL_ARM_BIGENDIAN          implies  is_substr(CYGBLD_GLOBAL_CFLAGS, " -mbig-endian ") }
        requires    { !CYGHWR_HAL_ARM_BIGENDIAN          implies !is_substr(CYGBLD_GLOBAL_CFLAGS, " -mbig-endian ") }
    }
    
    cdl_option CYGBLD_ARCH_LDFLAGS {
        display     "Architecture-specific linker flags"
        parent      CYGBLD_GLOBAL_OPTIONS
        flavor      data
        no_define
        calculated  { (CYGHWR_THUMB ? " -mthumb " : "") .
            (CYGBLD_ARM_ENABLE_THUMB_INTERWORK ? " -mthumb-interwork " : " -mno-thumb-interwork ") .
            (CYGHWR_HAL_ARM_BIGENDIAN ? " -mbig-endian " : "")
        }
        requires    {  CYGHWR_THUMB &&  CYGBLD_ARM_ENABLE_THUMB_INTERWORK implies  is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mthumb ") &&
                                                                                   is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mthumb-interwork ") &&
                                                                                  !is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mno-thumb-interwork ") }
        requires    { !CYGHWR_THUMB &&  CYGBLD_ARM_ENABLE_THUMB_INTERWORK implies !is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mthumb ") &&
                                                                                   is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mthumb-interwork ") &&
                                                                                  !is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mno-thumb-interwork ") }
        requires    {  CYGHWR_THUMB && !CYGBLD_ARM_ENABLE_THUMB_INTERWORK implies  is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mthumb ") &&
                                                                                  !is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mthumb-interwork ") &&
                                                                                   is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mno-thumb-interwork ") }
        requires    { !CYGHWR_THUMB && !CYGBLD_ARM_ENABLE_THUMB_INTERWORK implies !is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mthumb ") &&
                                                                                  !is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mthumb-interwork ") &&
                                                                                   is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mno-thumb-interwork ") }
        requires    {  CYGHWR_HAL_ARM_BIGENDIAN          implies  is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mbig-endian ") }
        requires    { !CYGHWR_HAL_ARM_BIGENDIAN          implies !is_substr(CYGBLD_GLOBAL_LDFLAGS, " -mbig-endian ") }
    }
    
    cdl_interface CYGINT_HAL_ARM_ARCH_ARM7 {
        display "The platform uses a processor with an ARM7 core"
    }

    cdl_interface CYGINT_HAL_ARM_ARCH_ARM9 {
        display "The platform uses a processor with an ARM9 core"
    }

    cdl_interface CYGINT_HAL_ARM_ARCH_ARM_CORTEXA9 {
        display "The platform uses a processor with an ARM Cortex-A9 multicore"
    }

    cdl_interface CYGINT_HAL_ARM_ARCH_STRONGARM {
        display "The platform uses a processor with a StrongARM core"
    }

    cdl_interface CYGINT_HAL_ARM_ARCH_XSCALE {
        display "The platform uses a processor with a XScale core"
    }

    cdl_option CYGHWR_HAL_ARM_CPU_FAMILY {
        display       "ARM CPU family"
        flavor        data
        legal_values  { (CYGINT_HAL_ARM_ARCH_ARM7 != 0) ? "ARM7" : ""
                        (CYGINT_HAL_ARM_ARCH_ARM9 != 0) ? "ARM9" : ""
                        (CYGINT_HAL_ARM_ARCH_STRONGARM != 0) ? "StrongARM" : ""
			(CYGINT_HAL_ARM_ARCH_ARM_CORTEXA9 != 0) ? "ARM Cortex-A9 MP" : ""
                        (CYGINT_HAL_ARM_ARCH_XSCALE != 0) ? "XScale" : ""
                        "" }
        default_value  { (CYGINT_HAL_ARM_ARCH_ARM7 != 0) ? "ARM7" : 
                         (CYGINT_HAL_ARM_ARCH_ARM9 != 0) ? "ARM9" : 
                         (CYGINT_HAL_ARM_ARCH_STRONGARM != 0) ? "StrongARM" :
			 (CYGINT_HAL_ARM_ARCH_ARM_CORTEXA9 != 0) ? "ARM Cortex-A9 MP" :	
                         (CYGINT_HAL_ARM_ARCH_XSCALE != 0) ? "XScale" :
                         "unknown" }
        no_define
        description   "
             It is possible to optimize code for different
             ARM CPU families. This option selects which CPU to
             optimize for on boards that support multiple CPU types."
    }

    cdl_option CYGBLD_HAL_ARM_EABI {
        display          "Build for ARM EABI"
        default_value    { (is_substr(CYGBLD_GLOBAL_COMMAND_PREFIX, "-eabi") && \
                            !is_substr(CYGBLD_GLOBAL_CFLAGS, "-mabi=apcs-gnu") && \
                            !is_substr(CYGBLD_GLOBAL_CFLAGS, "-mabi=atpcs")) || \
                           is_substr(CYGBLD_GLOBAL_CFLAGS, "-mabi=aapcs") }
        # The EABI uses a different C++ exception implementation to the standard
        # one and thus we indicate this to CYGPKG_LIBSTDCXX
        implements       CYGINT_LIBSTDCXX_NO_CXX_EXCEPTION_REG_FRAME_IMPL
        description "
            If using a toolchain which targets the ARM EABI (embedded application
            binary interface), this option should be enabled to provide altered
            semantics and differing linker section output."
    }

    cdl_option CYGHWR_HAL_ARM_DUMP_EXCEPTIONS {
        display          "Provide diagnostic dump for exceptions"
        requires         !CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
        default_value    0
        description      "
            Print messages about hardware exceptions, including
            raw exception frame dump and register contents."
    }

    cdl_option CYGIMP_HAL_PROCESS_ALL_EXCEPTIONS {
        display          "Process all exceptions with the eCos application"
        default_value    0
        description      "
           Normal RAM-based programs which do not include GDB stubs 
           defer processing of the illegal instruction exception to GDB.
           Setting this options allows the program to explicitly handle
           the illegal instruction exception itself.  Note: this will
           prevent the use of GDB to debug the application as breakpoints
           will no longer work."
    }

    cdl_option CYGHWR_HAL_ARM_ICE_THREAD_SUPPORT {
        display          "Support GDB thread operations via ICE/Multi-ICE"
        default_value    0
        requires         CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
        requires         CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
        requires         CYGDBG_KERNEL_DEBUG_GDB_THREAD_SUPPORT
        description      "
           Allow GDB to get thread information via the ICE/Multi-ICE
           connection."
    }

    cdl_option CYGOPT_HAL_ARM_SYSCALL_GPROF_SUPPORT {
	display		"Support for 'gprof' callbacks"
	calculated	1
	no_define
	active_if	CYGSEM_REDBOOT_BSP_SYSCALLS
	active_if	{ CYGDBG_HAL_DEBUG_GDB_CTRLC_SUPPORT || CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT }
	implements	CYGINT_REDBOOT_BSP_SYSCALLS_GPROF_SUPPORT
	description	"
	    The ARM HAL provides the macro for 'gprof' callbacks from RedBoot
	    to acquire the interrupt-context PC and SP, when this option is
            active."
    }

    cdl_option CYGOPT_HAL_ARM_WITH_USER_MODE {
        display          "Accept exceptions and irq's occurring in user mode"
        default_value    0
        description      "
            For standalone Redboot based programs running in user mode."
    }

    cdl_option CYGOPT_HAL_ARM_PRESERVE_SVC_SPSR {
        display          "Preserve svc spsr before returning to svc mode"
        default_value    0
        description      "
            This option secures exception and breakpoint processing
            triggered during execution of application specific SWI
            handlers."
    }

    cdl_option CYGOPT_HAL_ARM_FIQ_DISABLE {
        display          "Disable FIQs"
        default_value    1
        description      "This option causes the HAL to disable both IRQ and FIQ
                          interrupts during critical sections. Disabling this option
                          causes eCos to only disable IRQs and puts FIQ
                          interrupts outside the eCos world where they cannot interact
                          with eCos in any way. Disabling this option also enables
                          a set of macros, HAL_DISABLE|ENABLE|RESTORE|QUERY_FIQ,
                          that provide control over the delivery of FIQs.
                          The default is for this option to be enabled, which provides
                          backward compatibility with previous versions of the ARM HAL."
    }

    cdl_option CYGNUM_HAL_ARM_FIQ_STACK_SIZE {
        display          "FIQ stack size"
        active_if        !CYGOPT_HAL_ARM_FIQ_DISABLE
        flavor           data
        legal_values     32 to 0x80000000
        default_value    512
        description      "This option set the size of the stack used to handle FIQ
                          interrupts. It is only used if the HAL is not disabling
                          FIQs during critical sections. Otherwise FIQs are translated
                          into IRQs and delivered on the standard interrupt stack."
    }
    
    
    cdl_component CYGPKG_REDBOOT_ARM_OPTIONS {
        display       "Redboot for ARM options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        cdl_component CYGPKG_REDBOOT_ARM_LINUX_EXEC {
            display        "Provide the exec command in RedBoot"
            flavor         none
            parent         CYGPKG_REDBOOT_ARM_OPTIONS
            active_if      CYGBLD_BUILD_REDBOOT_WITH_EXEC
            description    "
                This option contains requirements for booting linux
                from RedBoot. The component is enabled/disabled from
                RedBoots CDL."
            compile -library=libextras.a redboot_linux_exec.c

            cdl_option CYGHWR_REDBOOT_LINUX_EXEC_X_SWITCH {
                display "Enable -x switch for exec command."
                flavor bool
                default_value 0
                description "
                    This option allows bi-endian platforms to launch kernels
                    built for an endianess different than the RedBoot endianess"
            }
 
            cdl_option CYGHWR_REDBOOT_ARM_LINUX_EXEC_ADDRESS {
                display       "Physical base address of linux kernel"
                flavor        data
                default_value CYGHWR_REDBOOT_ARM_LINUX_EXEC_ADDRESS_DEFAULT
                description   "
                    This is the physical address of the base of the 
                    Linux kernel image."
            }

            cdl_option CYGHWR_REDBOOT_ARM_LINUX_EXEC_ADDRESS_DEFAULT {
                display       "Default physical base address of linux kernel"
                flavor        data
                default_value 0x00008000
                no_define
                description   "
                    This is the physical address of the base of the 
                    Linux kernel image. This option gets set by the 
                    platform CDL."
            }

            cdl_option CYGHWR_REDBOOT_ARM_LINUX_TAGS_ADDRESS {
                display       "Base address of linux kernel parameter tags"
                flavor        data
                default_value 0x100
                description   "
                   This is the base address of the area of memory used to
                   pass parameters to the Linux kernel. This should be chosen
                   to avoid overlap with the kernel and any ramdisk image."
            }
        }

    }

    cdl_option CYGBLD_HAL_ARM_MCOUNT {
        display           "Support call-graph profiling"
        flavor            bool
        no_define
        active_if         CYGPKG_PROFILE_GPROF
        calculated        CYGPKG_PROFILE_CALLGRAPH
        requires          { CYGHWR_THUMB implies CYGBLD_ARM_ENABLE_THUMB_INTERWORK }
        compile           mcount.S
        description       "
            Calculate whether mcount functions should be built
            to support call-graph profiling."
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
        display "Linker script"
        flavor data
	no_define
        calculated  { "src/arm.ld" }
    }

    cdl_interface CYGINT_HAL_ARM_MEM_REAL_REGION_TOP {
        display  "Implementations of hal_arm_mem_real_region_top()"
    }
}

# EOF hal_arm.cdl
