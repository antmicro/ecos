# ====================================================================
#
#      wallclock_ds1307.cdl
#
#      eCos configuration data for Dallas 1307
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003, 2004 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:   jskov
# Date:           2001-07-06
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVICES_WALLCLOCK_DALLAS_DS1307 {
    parent        CYGPKG_IO_WALLCLOCK
    active_if     CYGPKG_IO_WALLCLOCK
    display       "Wallclock device driver for Dallas 1307"
    description   "
        This package provides a file with init, get and set functions
        for the Dallas 1307 clock part."
    doc           ref/devs-wallclock-dallas-ds1307-part.html

    compile       ds1307.cxx

    implements    CYGINT_WALLCLOCK_HW_IMPLEMENTATIONS
    active_if     CYGIMP_WALLCLOCK_HARDWARE
    implements    CYGINT_WALLCLOCK_SET_GET_MODE_SUPPORTED

    cdl_option CYGIMP_WALLCLOCK_HARDWARE {
        parent    CYGPKG_IO_WALLCLOCK_IMPLEMENTATION
        display       "Hardware wallclock"
        default_value 1
        implements    CYGINT_WALLCLOCK_IMPLEMENTATIONS
    }

    cdl_interface CYGINT_DEVICES_WALLCLOCK_DALLAS_DS1307_I2C {
	display		"Access DS1307 device via the I2C API"
	flavor		bool
	description "
            This interface will be implemented if the platform supports
            the standard I2C API and the platform HAL exports an I2C
            device cyg_i2c_wallclock_ds1307."
    }
    
    cdl_component CYGPKG_DEVICES_WALLCLOCK_DALLAS_DS1307_OPTIONS {
        display "DS1307 wallclock build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_DEVICES_WALLCLOCK_DALLAS_DS1307_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the wallclock device. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_DEVICES_WALLCLOCK_DALLAS_DS1307_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the wallclock device. These flags are removed from
                the set of global flags if present."
        }

    }
}
