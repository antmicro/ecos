##==========================================================================
##
##      hal_cortexm_stm32_stm3210e_eval.cdl
##
##      Cortex-M STM3210E EVAL platform HAL configuration data
##
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008, 2012 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##==========================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):    nickg
## Date:         2008-07-30
##
######DESCRIPTIONEND####
##
##==========================================================================

cdl_package CYGPKG_HAL_CORTEXM_STM32_STM3210E_EVAL {
    display       "ST STM3210E EVAL Development Board HAL"
    parent        CYGPKG_HAL_CORTEXM_STM32
    requires      { CYGHWR_HAL_CORTEXM_STM32_FAMILY == "F1" }
    requires      { CYGHWR_HAL_CORTEXM_STM32_F1 == "F103ZE" }
    define_header hal_cortexm_stm32_stm3210e_eval.h
    include_dir   cyg/hal
    hardware
    description   "
        The STM3210E EVAL HAL package provides the support needed to run
        eCos on the ST STM3210E EVAL board."

    compile       stm3210e_eval_misc.c

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_cortexm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_cortexm_stm32.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_cortexm_stm32_stm3210e_eval.h>"
	puts $::cdl_header "#define HAL_PLATFORM_CPU    \"Cortex-M3\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"ST STM3210E EVAL\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        default_value {"RAM"}
        legal_values  {"RAM" "SRAM" "ROM" "JTAG"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
            When targetting the ST STM3210E EVAL board it is possible to
            build the system for either RAM bootstrap or ROM bootstrap.
            Select 'RAM' when building programs to load into RAM using onboard
            debug software such as RedBoot or eCos GDB stubs.  Select 'ROM'
            when building a stand-alone application which will be put
            into ROM. The 'JTAG' type allows programs to be downloaded using a
            JTAG debugger such as a BDI3000 or PEEDI. The 'SRAM' type allows
            programs to be downloaded via a JTAG debugger into on-chip SRAM."
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated    { (CYG_HAL_STARTUP == "RAM" ) ? 
                        (CYGMEM_HAL_CORTEXM_STM32_STM3210E_EXTRA_BASE_RAM ?
                        "cortexm_stm3210e_eval_extrabaseram" : "cortexm_stm3210e_eval_ram")      :
                        (CYG_HAL_STARTUP == "SRAM") ? "cortexm_stm3210e_eval_sram"     :
                        (CYG_HAL_STARTUP == "ROM" ) ? "cortexm_stm3210e_eval_rom"      :
                        (CYG_HAL_STARTUP == "JTAG") ? "cortexm_stm3210e_eval_jtag"     :
                                                      "undefined" }

        cdl_option CYGMEM_HAL_CORTEXM_STM32_STM3210E_EXTRA_BASE_RAM {
            display       "Additional reserved space at base of RAM"
            flavor        booldata
            default_value 0
            active_if     {CYG_HAL_STARTUP == "RAM"}
            legal_values  0 to 0x80000
            description   "
                If you are using a RedBoot with additional components enabled,
                such as networking, RedBoot may be occupying additional RAM.
                In such cases, an eCos application loaded by RedBoot must
                reserve additional space at the base of RAM to accommodate
                RedBoot's extra RAM requirements. This option, specified in
                bytes, allows the amount of extra reserved space to be
                increased beyond the default."
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
                display "Memory layout linker script fragment"
                flavor data
                no_define
                define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
                calculated { "<pkgconf/mlt_" . CYGHWR_MEMORY_LAYOUT . ".ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
                display "Memory layout header file"
                flavor data
                no_define
                define -file system.h CYGHWR_MEMORY_LAYOUT_H
                calculated { "<pkgconf/mlt_" . CYGHWR_MEMORY_LAYOUT . ".h>" }
        }

    }

    cdl_option CYGARC_HAL_CORTEXM_STM32_INPUT_CLOCK {
        display         "Input Clock frequency"
        flavor          data
        default_value   8000000
        legal_values    0 to 1000000000
        description     "Main clock input."
    }

    cdl_component CYGHWR_HAL_CORTEXM_STM32_FLASH {
        display         "Flash support"
        parent          CYGPKG_IO_FLASH
        active_if       CYGPKG_IO_FLASH
        compile         -library=libextras.a stm3210e_eval_flash.c
        default_value   1
        description     "Control flash device support for STM3210E-EVAL board."
    
        cdl_option CYGHWR_HAL_CORTEXM_STM32_FLASH_INTERNAL {
            display         "Internal flash support"
            default_value   1
            description     "This option enables support for the internal flash device."
        }

        cdl_option CYGHWR_HAL_CORTEXM_STM32_FLASH_NOR {
            display         "External NOR flash support"
            default_value   1
            description     "This option enables support for the external NOR flash device."
        }

    }

    # Both UARTs 0 and 1 are available for diagnostic/debug use.
    implements CYGINT_HAL_STM32_UART0
    implements CYGINT_HAL_STM32_UART1

    implements      CYGINT_IO_SERIAL_FLOW_CONTROL_HW
    implements      CYGINT_IO_SERIAL_LINE_STATUS_HW
    
    
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   2
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The ST STM3210E EVAL board has two serial ports. This option
            chooses which port will be used to connect to a host
            running GDB."
     }

     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    0
         description      "
            The ST STM3210E EVAL has two serial ports. This option
            chooses which port will be used for diagnostic output."
     }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Console serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 38400
        description   "
            This option controls the default baud rate used for the
            console connection.
            RedBoot usess polling to transfer data over this port and
            might not be able to keep up with baud rates above the
            default, particularly when doing XYZmodem downloads. The
            interrupt-driven device driver is able to handle these
            baud rates, so any high speed application transfers should
            use that instead.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 38400
        description   "
            This option controls the default baud rate used for the
            GDB connection.
            RedBoot usess polling to transfer data over this port and
            might not be able to keep up with baud rates above the
            default, particularly when doing XYZmodem downloads. The
            interrupt-driven device driver is able to handle these
            baud rates, so any high speed application transfers should
            use that instead.
            Note: this should match the value chosen for the console port if the
            console and GDB port are the same."
    }

    cdl_component CYGHWR_HAL_CORTEXM_STM32_SPIETH_CONTROLLER {
        display       "STM3210E support for ENC424J600 SPI ethernet"
        parent        CYGPKG_DEVS_ETH_ENC424J600
        active_if     CYGPKG_DEVS_ETH_ENC424J600
        compile       stm3210e_eval_eth_enc424j600.c
        flavor        none
        no_define

        description   "
            Support for ENC424J600 with STM3210E EVAL board."
            
        cdl_option CYGNUM_ETH_SPIETH_HAL_INTERRUPT_VECTOR { 
            display       "Interrupt vector calculated from pin"
            parent        CYGNUM_DEVS_ETH_ENC424J600_INTERRUPT_VECTOR
            flavor        data
            no_define
            calculated    { "CYGNUM_HAL_INTERRUPT_EXTI" . CYGHWR_HAL_SPIETH_INTERRUPT_PIN } 
            active_if     CYGINT_IO_ETH_INT_SUPPORT_REQUIRED 
            description   "
                Interrupt vector corresponding with external interrupt line used for
                enc424j600.
                This value is automatically calculated from CYGHWR_HAL_SPIETH_INTERRUPT_PIN.
                "
        } 

        cdl_option CYGHWR_HAL_CORTEXM_STM32_SPIETH_SPI_BUS {
            display       "SPI bus"
            flavor        data
            requires      { (CYGHWR_HAL_CORTEXM_STM32_SPIETH_SPI_BUS == 1) implies CYGHWR_DEVS_SPI_CORTEXM_STM32_BUS1 }
            requires      { (CYGHWR_HAL_CORTEXM_STM32_SPIETH_SPI_BUS == 2) implies CYGHWR_DEVS_SPI_CORTEXM_STM32_BUS2 }
            requires      { (CYGHWR_HAL_CORTEXM_STM32_SPIETH_SPI_BUS == 3) implies CYGHWR_DEVS_SPI_CORTEXM_STM32_BUS3 }
            requires      (CYGNUM_DEVS_SPI_CORTEXM_STM32_PIN_TOGGLE_RATE==50)
            legal_values  { 1 2 3 } 
            default_value 1
            description   "
                Select which SPI bus of the STM32 the SPI Ethernet controller
                is connected to."
        }
        
        cdl_option CYGHWR_HAL_CORTEXM_STM32_SPIETH_SPI_CS {
            display       "Chip select index"
            flavor        data
            default_value 0
            legal_values  0 to 99
            description   "
                Enter the index into the array of chip selects to be used as
                the chip select for the external Ethernet
                controller connected to the SPI bus. The list of possible chip
                selects for the selected SPI bus is defined in the STM32 SPI
                driver's configuration, for example for SPI bus 1:
                CYGHWR_DEVS_SPI_CORTEXM_STM32_BUS1_CS_GPIOS."
        }
        
        cdl_option CYGHWR_HAL_CORTEXM_STM32_SPIETH_INTERRUPT_PORT {
            display       "Interrupt pin port"
            active_if     CYGINT_IO_ETH_INT_SUPPORT_REQUIRED 
            flavor        data
            legal_values  { "\'A\'" "\'B\'" "\'C\'" "\'D\'" "\'E\'" "\'F\'" "\'G\'" }
            default_value {"\'G\'"}
            description   "
               This selects the GPIO port associated with the interrupt pin
               connected to the external Ethernet controller."
        }
        
        cdl_option CYGHWR_HAL_SPIETH_INTERRUPT_PIN {
            display       "Interrupt pin number"
            active_if     CYGINT_IO_ETH_INT_SUPPORT_REQUIRED 
            flavor        data
            legal_values  0 to 15
            default_value 15
            description   "
               This selects the pin number within the GPIO port associated with
               the interrupt pin connected to the external Ethernet controller."
        }

        cdl_option CYGNUM_HAL_SPIETH_INTERRUPT_PRIORITY {
            display       "Interrupt priority"
            active_if     CYGINT_IO_ETH_INT_SUPPORT_REQUIRED 
            flavor        data
            legal_values  { 0xe0 0xd0 0xc0 0xb0 0xa0 0x90 0x80
                            0x70 0x60 0x50 0x40 0x30 0x20 0x10 0x00}
            default_value 0xe0
            description   "
               Enter the interrupt priority used for the interrupt
               connected to the external Ethernet controller. A
               lower number means a higher priority."
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-eabi" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGBLD_GLOBAL_WARNFLAGS . "-mcpu=cortex-m3 -mthumb -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-mcpu=cortex-m3 -mthumb -Wl,--gc-sections -Wl,-static -Wl,-n -g -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
    }

    cdl_component CYGPKG_HAL_CORTEXM_STM32_STM3210E_EVAL_OPTIONS {
        display "stm3210e HAL build options"
                flavor  none
                description   "
                        Package specific build options including control over
                        compiler flags used only in building this HAL."

                cdl_option CYGPKG_HAL_CORTEXM_STM32_STM3210E_EVAL_CFLAGS_ADD {
                        display "Additional compiler flags"
                        flavor  data
                        no_define
                        default_value { "-Werror" }
                        description   "
                                This option modifies the set of compiler flags
                                for building this HAL. These flags are used
                                in addition to the set of global flags."
                        }
                cdl_option CYGPKG_HAL_CORTEXM_STM32_STM3210E_EVAL_CFLAGS_REMOVE {
                        display "Suppressed compiler flags"
                        flavor  data
                        no_define
                        default_value { "" }
                        description   "
                                This option modifies the set of compiler flags
                                for building this HAL. These flags are
                                removed from the set of global flags if
                                present."
                }
        }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" || CYG_HAL_STARTUP == "JTAG" }
        requires      { CYGDBG_HAL_CRCTABLE_LOCATION == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "Generic" "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             Firstly there is \"Generic\" support which prevents the HAL
             from overriding the hardware vectors that it does not use, to
             instead allow an installed ROM monitor to handle them. This is
             the most basic support which is likely to be common to most
             implementations of ROM monitor.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
     }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        requires { CYGNUM_REDBOOT_FLASH_BASE == 0x64000000 }
        requires { CYGBLD_REDBOOT_MAX_MEM_SEGMENTS == 2 }

        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary images"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to binary image formats suitable for ROM programming."

            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img)
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

    cdl_component CYGBLD_HAL_CORTEXM_STM3210E_EVAL_GDB_STUBS {
        display "Create StubROM SREC and binary files"
        active_if CYGBLD_BUILD_COMMON_GDB_STUBS
        no_define
        calculated 1
        requires { CYG_HAL_STARTUP == "ROM" }

        make -priority 325 {
                <PREFIX>/bin/stubrom.srec : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O srec $< $@
        }
        make -priority 325 {
                <PREFIX>/bin/stubrom.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O binary $< $@
        }

        description "This component causes the ELF image generated by the
                     build process to be converted to S-Record and binary
                     files."
    }
}
