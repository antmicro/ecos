# ====================================================================
#
#      ser_mips_vrc437x.cdl
#
#      eCos serial MIPS/VRC437X configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  gthomas
# Contributors:
# Date:           1999-07-14
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_MIPS_VRC437X {
    display       "VRC437X serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_MIPS_VR4300_VRC437X

    requires      CYGPKG_ERROR
    include_dir   cyg/io
    include_files ; # none _exported_ whatsoever
    description   "
           This option enables the serial device drivers for the
           VRC437X."

    compile       -library=libextras.a   vrc437x_serial.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_mips_vrc437x.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

cdl_component CYGPKG_IO_SERIAL_MIPS_VRC437X_SERIAL0 {
    display       "VRC437X serial port 0 driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for the VRC437X port 0."

    cdl_option CYGDAT_IO_SERIAL_MIPS_VRC437X_SERIAL0_NAME {
        display       "Device name for the VRC437X serial port 0 driver"
        flavor        data
        default_value {"\"/dev/ser0\""}
        description   "
            This option sets the name of the serial device for the VRC437X 
            port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_MIPS_VRC437X_SERIAL0_BAUD {
        display       "Baud rate for the VRC437X serial port 0 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
            VRC437X port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_MIPS_VRC437X_SERIAL0_BUFSIZE {
        display       "Buffer size for the VRC437X serial port 0 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used
            for the VRC437X port 0."
    }
}
cdl_component CYGPKG_IO_SERIAL_MIPS_VRC437X_SERIAL1 {
    display       "VRC437X serial port 1 driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for the VRC437X port 1."

    cdl_option CYGDAT_IO_SERIAL_MIPS_VRC437X_SERIAL1_NAME {
        display       "Device name for the VRC437X serial port 1 driver"
        flavor        data
        default_value {"\"/dev/ser1\""}
        description   "
            This option specifies the name of serial device for the
            VRC437X port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_MIPS_VRC437X_SERIAL1_BAUD {
        display       "Baud rate for the VRC437X serial port 1 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
            VRC437X port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_MIPS_VRC437X_SERIAL1_BUFSIZE {
        display       "Buffer size for the VRC437X serial port 1 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used for
            the VRC437X port 1."
    }
}

    cdl_component CYGPKG_IO_SERIAL_MIPS_VRC437X_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_MIPS_VRC437X_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_MIPS_VRC437X_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_MIPS_VRC437X_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_IO_SERIAL_MIPS_VRC437X_SERIAL0

        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_MIPS_VRC437X_SERIAL0_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"vrc437X\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty0\""
        }
    }
}

# EOF ser_mips_vrc437x.cdl
