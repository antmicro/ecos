# ====================================================================
#
#      ser_arm_at91.cdl
#
#      eCos serial Atmel AT91 (ARM) configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Contributors:   tkoeller
# Date:           2001-07-24
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_ARM_AT91 {
    display       "Atmel AT91 serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_ARM_AT91

    requires      CYGPKG_ERROR
    include_dir   cyg/io
    include_files ; # none _exported_ whatsoever
    description   "
           This option enables the serial device drivers for the
           Atmel AT91."
    
    implements    CYGINT_IO_SERIAL_BLOCK_TRANSFER

    compile       -library=libextras.a   at91_serial.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_arm_at91.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

cdl_component CYGPKG_IO_SERIAL_ARM_AT91_SERIAL0 {
    display       "Atmel AT91 serial port 0 driver"
    flavor        bool
    default_value 0
    description   "
        This option includes the serial device driver for the Atmel AT91 
        port 0 (serial A)."

    cdl_option CYGDAT_IO_SERIAL_ARM_AT91_SERIAL0_NAME {
        display       "Device name for Atmel AT91 serial port 0 driver"
        flavor        data
        default_value {"\"/dev/ser0\""}
        description   "
            This option specifies the name of the serial device for the 
            Atmel AT91 port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_ARM_AT91_SERIAL0_BAUD {
        display       "Baud rate for the Atmel AT91 serial port 0 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the 
            Atmel AT91 port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_ARM_AT91_SERIAL0_BUFSIZE {
        display       "Buffer size for the Atmel AT91 serial port 0 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the Atmel AT91 port 0."
    }
    
    cdl_option CYGNUM_IO_SERIAL_ARM_AT91_SERIAL0_RCV_CHUNK_SIZE {
        display       "Receive data chunk size"
        flavor        data
        legal_values  1 to 65519
        default_value 1
        description   "
            This parameter can be used to reduce the number of interrupts
            that must be processed by the driver. An interrupt will only
            be generated if either this many data bytes have been received
            or the receiver has been idle for some time. This reduces
            overall system load at the expense of making the driver less
            responsive and using slightly more memory for buffering data.
            Setting this parameter to 1 will give standard behavior."
    }
}

cdl_component CYGPKG_IO_SERIAL_ARM_AT91_SERIAL1 {
    display       "Atmel AT91 serial port 1 driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for the Atmel AT91 
        port 1 (serial B)."

    cdl_option CYGDAT_IO_SERIAL_ARM_AT91_SERIAL1_NAME {
        display       "Device name for Atmel AT91 serial port 1 driver"
        flavor        data
        default_value {"\"/dev/ser1\""}
        description   "
            This option specifies the name of the serial device for the 
            Atmel AT91 port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_ARM_AT91_SERIAL1_BAUD {
        display       "Baud rate for the Atmel AT91 serial port 1 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
            Atmel AT91 port 1."
    }

    cdl_option CYGNUM_IO_SERIAL_ARM_AT91_SERIAL1_BUFSIZE {
        display       "Buffer size for the Atmel AT91 serial port 1 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the Atmel AT91 port 1."
    }
    
    cdl_option CYGNUM_IO_SERIAL_ARM_AT91_SERIAL1_RCV_CHUNK_SIZE {
        display       "Receive data chunk size"
        flavor        data
        legal_values  1 to 65519
        default_value 1
        description   "
            This parameter can be used to reduce the number of interrupts
            that must be processed by the driver. An interrupt will only
            be generated if either this many data bytes have been received
            or the receiver has been idle for some time. This reduces
            overall system load at the expense of making the driver less
            responsive and using slightly more memory for buffering data.
            Setting this parameter to 1 will give standard behavior."
    }
}

cdl_component CYGPKG_IO_SERIAL_ARM_AT91_SERIAL2 {
    display       "Atmel AT91 serial port 2 driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for the Atmel AT91 
        port 2 (serial C)."

    cdl_option CYGDAT_IO_SERIAL_ARM_AT91_SERIAL2_NAME {
        display       "Device name for Atmel AT91 serial port 1 driver"
        flavor        data
        default_value {"\"/dev/ser2\""}
        description   "
            This option specifies the name of the serial device for the 
            Atmel AT91 port 2."
    }

    cdl_option CYGNUM_IO_SERIAL_ARM_AT91_SERIAL2_BAUD {
        display       "Baud rate for the Atmel AT91 serial port 1 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
            Atmel AT91 port 2."
    }

    cdl_option CYGNUM_IO_SERIAL_ARM_AT91_SERIAL2_BUFSIZE {
        display       "Buffer size for the Atmel AT91 serial port 2 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the Atmel AT91 port 2."
    }
    
    cdl_option CYGNUM_IO_SERIAL_ARM_AT91_SERIAL2_RCV_CHUNK_SIZE {
        display       "Receive data chunk size"
        flavor        data
        legal_values  1 to 65519
        default_value 1
        description   "
            This parameter can be used to reduce the number of interrupts
            that must be processed by the driver. An interrupt will only
            be generated if either this many data bytes have been received
            or the receiver has been idle for some time. This reduces
            overall system load at the expense of making the driver less
            responsive and using slightly more memory for buffering data.
            Setting this parameter to 1 will give standard behavior."
    }
}


    cdl_component CYGPKG_IO_SERIAL_ARM_AT91_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_ARM_AT91_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_ARM_AT91_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_AT91_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_IO_SERIAL_ARM_AT91_SERIAL1

        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_ARM_AT91_SERIAL1_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"eb40\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty1\""
        }
    }
}

# EOF ser_arm_at91.cdl
