#==========================================================================
# 
#       qspi_xc7z.cdl
# 
#       Xilinx XC7Z020 (ARM) QSPI driver configuration data
# 
#==========================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
#==========================================================================
######DESCRIPTIONBEGIN####
# 
# Author(s):    ITR GmbH
# Date:         2012-07-09
# Purpose:      
# Description:  QSPI driver for Xilinx XC7Z020 ARM Cortex-A9
# 
#####DESCRIPTIONEND####
# 
#==========================================================================

cdl_package CYGPKG_DEVS_QSPI_ARM_XC7Z {
    parent        CYGPKG_IO_SPI
    active_if     CYGPKG_IO_SPI
    display       "Xilinx XC7Z QSPI driver"
    requires      CYGPKG_HAL_ARM_XC7Z
    requires      CYGPKG_ERROR
    hardware
    include_dir   cyg/io
    compile       qspi_xc7z.c
    compile       -library=libextras.a qspi_xc7z_init.cxx

    cdl_option CYGHWR_DEVS_QSPI_ARM_XC7Z {
        display       "Enable support for QSPI"
        flavor        bool
        default_value 1
        description   "Enable this option to add support for the first 
                QSPI peripheral. The most XC7Z devices only have one bus" 
    }

    cdl_component CYGPKG_DEVS_QSPI_ARM_XC7Z_OPTIONS {
        display "Xilinx XC7Z QSPI driver build options"
        flavor  none
        description   "
            Package specific build options including control over
            compiler flags used only in building this package,
            and details of which tests are built."

        cdl_option CYGPKG_DEVS_QSPI_ARM_XC7Z_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the QSPI device. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_DEVS_QSPI_ARM_XC7Z_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the QSPI device. These flags are removed from
                the set of global flags if present."
        }
    }
}

# EOF qspi_xc7z.cdl